magic
tech scmos
timestamp 1543950581
<< metal1 >>
rect -24 174 219 177
rect -24 168 -1 174
rect 64 168 69 174
rect 213 168 219 174
rect 31 96 35 109
rect -24 78 -1 96
rect 64 83 219 96
rect 64 78 87 83
rect 93 78 219 83
rect 1 53 5 78
rect 193 58 219 62
rect 86 54 87 58
rect 66 48 68 52
rect -2 42 -1 46
rect 67 38 71 42
rect -10 24 8 28
rect -17 17 8 21
rect -24 1 87 6
rect 93 1 219 6
rect -24 -3 219 1
<< m2contact >>
rect 23 128 27 132
rect 15 105 19 109
rect 189 58 193 62
rect 68 48 72 52
rect -6 42 -2 46
rect 61 38 65 42
rect -14 24 -10 28
rect 8 24 12 28
rect -21 17 -17 21
rect 8 17 12 21
<< metal2 >>
rect -21 21 -17 177
rect -21 -3 -17 17
rect -14 28 -10 177
rect 1 164 5 177
rect 152 173 156 177
rect 204 142 208 171
rect 27 128 49 132
rect 160 130 213 134
rect 45 116 49 128
rect 65 119 69 123
rect 19 106 49 109
rect 19 105 35 106
rect 45 89 49 106
rect 45 85 193 89
rect 58 71 87 75
rect 189 62 193 85
rect -14 -3 -10 24
rect -6 10 -2 42
rect 12 24 56 28
rect 61 24 65 38
rect 68 21 72 48
rect 12 17 56 21
rect 62 17 72 21
rect 1 -3 5 10
rect 208 4 212 86
rect 152 0 212 4
rect 152 -3 156 0
<< m3contact >>
rect 203 171 208 176
rect 213 129 218 134
rect -7 5 -2 10
<< metal3 >>
rect 202 176 209 177
rect 202 171 203 176
rect 208 171 209 176
rect 202 170 209 171
rect 212 134 219 135
rect 212 129 213 134
rect 218 129 219 134
rect 212 95 219 129
rect -8 10 209 11
rect -8 5 -7 10
rect -2 5 209 10
rect -8 4 209 5
rect 202 -3 209 4
use ../../fa/magic/fa  fa_0 ../../fa/magic
timestamp 1543290821
transform 1 0 39 0 1 90
box 0 -4 175 87
use ../../bc1a/magic/bc1a  bc1a_0 ../../bc1a/magic
timestamp 1543295583
transform 1 0 0 0 1 12
box -1 -12 64 162
use ../../nand/magic/nand  nand_0 ../../nand/magic
timestamp 1543290081
transform 1 0 59 0 -1 81
box -4 -3 28 81
use ../../dffpos/magic/dffpos  dffpos_0 ../../dffpos/magic
timestamp 1543271063
transform 1 0 57 0 1 0
box 18 0 139 84
<< labels >>
rlabel metal2 154 175 154 175 0 Cin
rlabel metal2 154 -2 154 -2 0 Cout
rlabel metal2 3 0 3 0 1 Init
rlabel metal3 217 98 217 98 7 fa_in
rlabel space 7 51 7 51 1 muxB_in
rlabel space 16 104 16 104 1 reg_in
rlabel metal2 -12 -1 -12 -1 1 clk
rlabel metal2 -20 -1 -20 -1 2 en
rlabel metal1 -22 87 -22 87 3 gnd
rlabel metal1 -22 173 -22 173 5 vdd
rlabel metal1 -22 1 -22 1 1 vdd
rlabel metal1 217 60 217 60 7 Out
rlabel metal3 205 0 205 0 1 muxA_in
rlabel m3contact 205 175 205 175 5 add_out
<< end >>
