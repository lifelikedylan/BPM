magic
tech scmos
timestamp 1541616290
<< nwell >>
rect -5 64 124 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
rect 23 6 25 16
rect 31 6 33 16
rect 36 6 38 16
rect 44 6 46 16
rect 52 6 54 16
rect 60 6 62 16
rect 68 6 70 16
rect 77 6 79 16
rect 82 6 84 16
rect 87 6 89 16
rect 95 6 97 16
rect 111 6 113 16
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
rect 31 74 33 94
rect 36 74 38 94
rect 44 74 46 94
rect 52 74 54 94
rect 60 74 62 94
rect 68 74 70 94
rect 77 74 79 94
rect 82 74 84 94
rect 87 74 89 94
rect 95 74 97 94
rect 111 74 113 94
<< ndiffusion >>
rect 6 6 7 16
rect 9 6 10 16
rect 14 6 15 16
rect 17 6 18 16
rect 22 6 23 16
rect 25 6 26 16
rect 30 6 31 16
rect 33 6 36 16
rect 38 6 39 16
rect 43 6 44 16
rect 46 6 47 16
rect 51 6 52 16
rect 54 6 55 16
rect 59 6 60 16
rect 62 6 63 16
rect 67 6 68 16
rect 70 6 71 16
rect 76 6 77 16
rect 79 6 82 16
rect 84 6 87 16
rect 89 6 90 16
rect 94 6 95 16
rect 97 6 98 16
rect 110 6 111 16
rect 113 6 114 16
<< pdiffusion >>
rect 6 74 7 94
rect 9 74 10 94
rect 14 74 15 94
rect 17 74 18 94
rect 22 74 23 94
rect 25 74 26 94
rect 30 74 31 94
rect 33 74 36 94
rect 38 74 39 94
rect 43 74 44 94
rect 46 74 47 94
rect 51 74 52 94
rect 54 74 55 94
rect 59 74 60 94
rect 62 74 63 94
rect 67 74 68 94
rect 70 74 71 94
rect 76 74 77 94
rect 79 74 82 94
rect 84 74 87 94
rect 89 74 90 94
rect 94 74 95 94
rect 97 74 98 94
rect 110 74 111 94
rect 113 74 114 94
<< ndcontact >>
rect 2 6 6 16
rect 10 6 14 16
rect 18 6 22 16
rect 26 6 30 16
rect 39 6 43 16
rect 47 6 51 16
rect 55 6 59 16
rect 63 6 67 16
rect 71 6 76 16
rect 90 6 94 16
rect 98 6 102 16
rect 106 6 110 16
rect 114 6 118 16
<< pdcontact >>
rect 2 74 6 94
rect 10 74 14 94
rect 18 74 22 94
rect 26 74 30 94
rect 39 74 43 94
rect 47 74 51 94
rect 55 74 59 94
rect 63 74 67 94
rect 71 74 76 94
rect 90 74 94 94
rect 98 74 102 94
rect 106 74 110 94
rect 114 74 118 94
<< psubstratepcontact >>
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
rect 94 -2 98 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
rect 94 98 98 102
rect 110 98 114 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 36 94 38 96
rect 44 94 46 96
rect 52 94 54 96
rect 60 94 62 96
rect 68 94 70 96
rect 77 94 79 96
rect 82 94 84 96
rect 87 94 89 96
rect 95 94 97 96
rect 111 94 113 96
rect 7 37 9 74
rect 15 47 17 74
rect 23 57 25 74
rect 7 16 9 33
rect 15 16 17 43
rect 23 16 25 53
rect 31 48 33 74
rect 36 73 38 74
rect 44 73 46 74
rect 36 71 46 73
rect 31 16 33 44
rect 44 37 46 71
rect 52 47 54 74
rect 60 57 62 74
rect 68 65 70 74
rect 44 19 46 33
rect 36 17 46 19
rect 36 16 38 17
rect 44 16 46 17
rect 52 16 54 43
rect 60 16 62 53
rect 68 29 70 61
rect 77 57 79 74
rect 78 53 79 57
rect 75 31 77 53
rect 82 48 84 74
rect 87 56 89 74
rect 87 54 92 56
rect 75 29 79 31
rect 68 16 70 25
rect 77 16 79 29
rect 82 16 84 44
rect 90 37 92 54
rect 95 43 97 74
rect 111 64 113 74
rect 107 62 113 64
rect 95 41 99 43
rect 87 33 88 37
rect 87 16 89 33
rect 97 29 99 41
rect 95 27 99 29
rect 95 23 97 27
rect 107 26 113 29
rect 95 16 97 19
rect 111 16 113 26
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
rect 36 4 38 6
rect 44 4 46 6
rect 52 4 54 6
rect 60 4 62 6
rect 68 4 70 6
rect 77 4 79 6
rect 82 4 84 6
rect 87 4 89 6
rect 95 4 97 6
rect 111 4 113 6
<< polycontact >>
rect 23 53 27 57
rect 15 43 19 47
rect 7 33 11 37
rect 31 44 35 48
rect 67 61 71 65
rect 59 53 63 57
rect 51 43 55 47
rect 43 33 47 37
rect 74 53 78 57
rect 81 44 85 48
rect 67 25 71 29
rect 103 62 107 66
rect 88 33 92 37
rect 103 26 107 30
rect 93 19 97 23
<< metal1 >>
rect -5 102 122 103
rect -5 98 -2 102
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 62 102
rect 66 98 78 102
rect 82 98 94 102
rect 98 98 110 102
rect 114 98 122 102
rect -5 97 122 98
rect 10 94 14 97
rect 39 94 43 97
rect 55 94 59 97
rect 90 94 94 97
rect 106 94 110 97
rect 76 74 78 77
rect 3 71 6 74
rect 18 71 21 74
rect 3 68 21 71
rect 48 71 51 74
rect 63 71 66 74
rect 48 68 66 71
rect 30 62 67 65
rect 71 62 103 65
rect 22 53 23 57
rect 27 54 59 57
rect 63 54 74 57
rect 10 43 15 47
rect 19 44 31 47
rect 35 44 51 47
rect 55 44 81 47
rect 102 43 122 47
rect 2 33 7 37
rect 11 33 43 36
rect 47 33 88 36
rect 30 26 67 29
rect 71 26 103 29
rect 3 19 21 22
rect 3 16 6 19
rect 18 16 21 19
rect 48 19 66 22
rect 75 20 93 23
rect 48 16 51 19
rect 63 16 66 19
rect 73 16 74 20
rect 100 16 103 19
rect 102 13 103 16
rect 10 3 14 6
rect 39 3 43 6
rect 55 3 59 6
rect 90 3 94 6
rect 106 3 110 6
rect -5 2 122 3
rect -5 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 62 2
rect 66 -2 78 2
rect 82 -2 94 2
rect 98 -2 122 2
rect -5 -3 122 -2
<< m2contact >>
rect 26 70 30 74
rect 74 70 78 74
rect 98 70 102 74
rect 114 70 118 74
rect 26 62 30 66
rect 18 53 22 57
rect 98 43 102 47
rect 114 33 118 37
rect 26 25 30 29
rect 26 16 30 20
rect 74 16 78 20
rect 100 19 104 23
rect 114 16 118 20
<< metal2 >>
rect 74 74 78 77
rect 26 66 30 70
rect 27 29 30 62
rect 26 20 30 25
rect 74 20 78 70
rect 99 47 102 70
rect 99 23 102 43
rect 115 37 118 70
rect 99 19 100 23
rect 115 20 118 33
<< labels >>
rlabel nsubstratencontact 0 100 0 100 4 vdd
rlabel metal1 4 0 4 0 1 gnd
rlabel metal1 4 35 4 35 1 A
rlabel m2contact 116 35 116 35 1 Cout
rlabel metal1 12 45 12 45 1 B
rlabel m2contact 20 55 20 55 1 C
rlabel metal1 109 45 109 45 1 SUm
<< end >>
