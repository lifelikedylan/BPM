magic
tech scmos
timestamp 1543875729
<< metal1 >>
rect 10 1434 14 1438
rect 17 1408 21 1412
rect 277 1391 281 1395
rect 277 1384 281 1388
rect 17 1362 21 1366
rect 277 1362 281 1366
rect 277 1341 281 1359
rect 17 1316 21 1341
rect 498 1333 504 1337
rect 498 1325 504 1329
rect 277 1312 281 1316
rect 17 1305 21 1309
rect 232 1306 236 1310
rect 277 1305 281 1309
rect 498 1305 504 1310
rect 17 1228 21 1232
rect 277 1211 281 1215
rect 277 1204 281 1208
rect 17 1182 21 1186
rect 277 1182 281 1186
rect 277 1161 281 1179
rect 17 1136 21 1161
rect 498 1153 504 1157
rect 498 1145 504 1149
rect 277 1132 281 1136
rect 17 1125 21 1129
rect 232 1126 236 1130
rect 277 1125 281 1129
rect 498 1125 504 1130
rect 17 1048 21 1052
rect 277 1031 281 1035
rect 277 1024 281 1028
rect 17 1002 21 1006
rect 277 1002 281 1006
rect 277 981 281 999
rect 17 956 21 981
rect 498 973 504 977
rect 498 965 504 969
rect 277 952 281 956
rect 17 945 21 949
rect 232 946 236 950
rect 277 945 281 949
rect 498 945 504 950
rect 17 868 21 872
rect 277 851 281 855
rect 277 844 281 848
rect 17 822 21 826
rect 277 822 281 826
rect 277 801 281 819
rect 17 776 21 801
rect 498 793 504 797
rect 498 785 504 789
rect 277 772 281 776
rect 17 765 21 769
rect 232 766 236 770
rect 277 765 281 769
rect 498 765 504 770
rect 17 688 21 692
rect 277 671 281 675
rect 277 664 281 668
rect 17 642 21 646
rect 277 642 281 646
rect 277 621 281 639
rect 17 596 21 621
rect 498 613 504 617
rect 498 605 504 609
rect 277 592 281 596
rect 17 585 21 589
rect 232 586 236 590
rect 277 585 281 589
rect 498 585 504 590
rect 17 508 21 512
rect 277 491 281 495
rect 277 484 281 488
rect 17 462 21 466
rect 277 462 281 466
rect 277 441 281 459
rect 17 416 21 441
rect 498 433 504 437
rect 498 425 504 429
rect 277 412 281 416
rect 17 405 21 409
rect 232 406 236 410
rect 277 405 281 409
rect 498 405 504 410
rect 17 328 21 332
rect 277 311 281 315
rect 277 304 281 308
rect 17 282 21 286
rect 277 282 281 286
rect 17 236 21 261
rect 498 253 504 257
rect 498 245 504 249
rect 277 232 281 236
rect 17 225 21 229
rect 232 226 236 230
rect 277 225 281 229
rect 498 225 504 230
rect 17 148 21 152
rect 277 138 281 142
rect 277 131 281 135
rect 277 124 281 128
rect 17 102 21 106
rect 277 102 281 106
rect 17 56 21 81
rect 500 73 504 77
rect 500 65 504 69
rect 277 52 281 56
rect 17 45 21 49
rect 232 46 236 50
rect 277 45 281 49
rect 499 45 504 50
rect 0 -4 268 -3
rect 0 -8 3 -4
rect 7 -8 263 -4
rect 267 -8 268 -4
rect 0 -9 268 -8
rect 0 -13 275 -12
rect 0 -17 10 -13
rect 14 -17 270 -13
rect 274 -17 275 -13
rect 0 -18 275 -17
rect 0 -22 261 -21
rect 0 -26 256 -22
rect 260 -26 261 -22
rect 0 -27 261 -26
rect 0 -31 254 -30
rect 0 -35 249 -31
rect 253 -35 254 -31
rect 0 -36 254 -35
rect 0 -40 296 -39
rect 0 -44 32 -40
rect 36 -44 291 -40
rect 295 -44 296 -40
rect 0 -45 296 -44
<< m2contact >>
rect 284 1398 288 1402
rect 284 1218 288 1222
rect 284 1038 288 1042
rect 284 858 288 862
rect 284 678 288 682
rect 284 498 288 502
rect 284 318 288 322
rect 284 138 288 142
rect 249 3 253 7
rect 3 -8 7 -4
rect 263 -8 267 -4
rect 10 -17 14 -13
rect 270 -17 274 -13
rect 256 -26 260 -22
rect 249 -35 253 -31
rect 32 -44 36 -40
rect 291 -44 295 -40
<< metal2 >>
rect 183 1439 260 1443
rect 241 1401 245 1405
rect 3 -4 7 1284
rect 10 -13 14 1291
rect 32 -40 36 1273
rect 241 1221 245 1225
rect 241 1041 245 1045
rect 241 861 245 865
rect 241 681 245 685
rect 241 501 245 505
rect 241 321 245 325
rect 241 141 245 145
rect 249 7 253 1436
rect 183 0 187 3
rect 249 -31 253 3
rect 256 -22 260 1439
rect 263 -4 267 1284
rect 270 -13 274 1291
rect 284 1222 288 1398
rect 284 1042 288 1218
rect 284 862 288 1038
rect 284 682 288 858
rect 284 502 288 678
rect 284 322 288 498
rect 284 142 288 318
rect 291 -40 295 1273
use ../../bs1/magic/bs1  bs1_0 ../../bs1/magic
array 0 0 245 0 7 180
timestamp 1543618603
transform 1 0 31 0 1 3
box -31 -3 214 177
use ../../bs2/magic/bs2  bs2_0 ../../bs2/magic
array 0 0 257 0 7 180
timestamp 1543628271
transform 1 0 290 0 1 3
box -46 -3 214 177
<< labels >>
rlabel metal1 2 -15 2 -15 2 clk
rlabel metal1 2 -6 2 -6 3 en
rlabel metal1 2 -33 2 -33 2 vdd
rlabel metal1 2 -24 2 -24 3 gnd
rlabel metal1 2 -42 2 -42 2 init
rlabel metal1 19 104 19 104 1 q_15
rlabel metal1 19 284 19 284 1 q_14
rlabel metal1 19 464 19 464 1 q_13
rlabel metal1 19 644 19 644 1 q_12
rlabel metal1 19 824 19 824 1 q_11
rlabel metal1 19 1004 19 1004 1 q_10
rlabel metal1 19 1184 19 1184 1 q_9
rlabel metal1 19 1364 19 1364 1 q_8
rlabel metal1 234 48 234 48 1 q_15
rlabel metal1 234 228 234 228 1 q_14
rlabel metal1 234 408 234 408 1 q_13
rlabel metal1 234 588 234 588 1 q_12
rlabel metal1 234 768 234 768 1 q_11
rlabel metal1 234 948 234 948 1 q_10
rlabel metal1 233 1128 233 1128 1 q_9
rlabel metal1 279 104 279 104 1 q_7
rlabel metal1 279 126 279 126 1 mplier_7
rlabel metal1 279 133 279 133 1 mcand_7
rlabel metal1 279 284 279 284 1 q_6
rlabel metal1 279 306 279 306 1 mplier_6
rlabel metal1 279 313 279 313 1 mcand_6
rlabel metal1 279 464 279 464 1 q_5
rlabel metal1 279 486 279 486 1 mplier_5
rlabel metal1 279 493 279 493 1 mcand_5
rlabel metal1 279 644 279 644 1 q_4
rlabel metal1 279 666 279 666 1 mplier_4
rlabel metal1 279 673 279 673 1 mcand_4
rlabel metal1 279 824 279 824 1 q_3
rlabel metal1 279 846 279 846 1 mplier_3
rlabel metal1 279 853 279 853 1 mcand_3
rlabel metal1 279 1004 279 1004 1 q_2
rlabel metal1 279 1026 279 1026 1 mplier_2
rlabel metal1 279 1033 279 1033 1 mcand_2
rlabel metal1 279 1184 279 1184 1 q_1
rlabel metal1 279 1206 279 1206 1 mplier_1
rlabel metal1 279 1213 279 1213 1 mcand_1
rlabel metal1 279 1386 279 1386 1 mplier_0
rlabel metal1 279 1393 279 1393 1 mcand_0
rlabel metal1 502 47 502 47 7 q_7
rlabel metal1 502 227 502 227 7 q_6
rlabel metal1 502 407 502 407 7 q_5
rlabel metal1 502 587 502 587 7 q_4
rlabel metal1 502 767 502 767 7 q_3
rlabel metal1 502 947 502 947 7 q_2
rlabel metal1 502 1128 502 1128 7 q_1
rlabel metal1 502 1307 502 1307 7 q_0
rlabel metal2 185 1 185 1 1 cout
rlabel metal1 234 1308 234 1308 1 q_8
<< end >>
