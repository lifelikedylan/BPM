magic
tech scmos
timestamp 1542251572
<< metal1 >>
rect -1 174 244 177
rect 64 168 69 174
rect 236 168 244 174
rect -1 145 8 149
rect 64 78 244 96
rect -1 -3 244 6
<< m2contact >>
rect 8 145 12 149
<< metal2 >>
rect 12 145 79 149
rect 75 123 79 145
rect 75 119 88 123
rect 60 112 67 116
rect 60 102 64 112
use ../../fa/magic/fa  fa_0 ../../fa/magic
timestamp 1542251572
transform 1 0 61 0 1 90
box 0 -4 175 89
use ../../bc1a/magic/bc1a  bc1a_0 ../../bc1a/magic
timestamp 1542169151
transform 1 0 0 0 1 12
box -1 -12 64 162
<< labels >>
rlabel metal1 176 176 176 176 5 c_in
rlabel metal1 1 147 1 147 3 fa_in
<< end >>
