magic
tech scmos
timestamp 1543271063
<< ntransistor >>
rect 33 65 35 75
rect 38 65 40 75
rect 54 65 56 75
rect 59 65 61 75
rect 67 65 69 75
rect 72 65 74 75
rect 81 65 83 75
rect 97 65 99 75
rect 102 65 104 75
rect 110 65 112 75
rect 115 65 117 75
rect 124 65 126 75
rect 129 65 131 75
<< ptransistor >>
rect 33 9 35 29
rect 38 9 40 29
rect 54 9 56 29
rect 59 9 61 29
rect 67 9 69 29
rect 72 9 74 29
rect 81 9 83 29
rect 97 9 99 29
rect 102 9 104 29
rect 110 9 112 29
rect 115 9 117 29
rect 124 9 126 29
rect 129 9 131 29
<< ndiffusion >>
rect 32 65 33 75
rect 35 65 38 75
rect 40 65 41 75
rect 53 65 54 75
rect 56 65 59 75
rect 61 65 62 75
rect 66 65 67 75
rect 69 65 72 75
rect 74 65 75 75
rect 80 65 81 75
rect 83 65 84 75
rect 96 65 97 75
rect 99 65 102 75
rect 104 65 105 75
rect 109 65 110 75
rect 112 65 115 75
rect 117 65 118 75
rect 123 65 124 75
rect 126 65 129 75
rect 131 65 132 75
<< pdiffusion >>
rect 32 9 33 29
rect 35 9 38 29
rect 40 9 41 29
rect 53 9 54 29
rect 56 9 59 29
rect 61 9 62 29
rect 66 9 67 29
rect 69 9 72 29
rect 74 9 75 29
rect 80 9 81 29
rect 83 9 84 29
rect 96 9 97 29
rect 99 9 102 29
rect 104 9 105 29
rect 109 9 110 29
rect 112 9 115 29
rect 117 9 118 29
rect 123 9 124 29
rect 126 9 129 29
rect 131 9 132 29
<< ndcontact >>
rect 28 65 32 75
rect 41 65 45 75
rect 49 65 53 75
rect 62 65 66 75
rect 75 65 80 75
rect 84 65 88 75
rect 92 65 96 75
rect 105 65 109 75
rect 118 65 123 75
rect 132 65 136 75
<< pdcontact >>
rect 28 9 32 29
rect 41 9 45 29
rect 49 9 53 29
rect 62 9 66 29
rect 75 9 80 29
rect 84 9 88 29
rect 92 9 96 29
rect 105 9 109 29
rect 118 9 123 29
rect 132 9 136 29
<< psubstratepcontact >>
rect 29 79 33 83
rect 37 79 41 83
rect 45 79 49 83
rect 53 79 57 83
rect 61 79 65 83
rect 69 79 73 83
rect 77 79 81 83
rect 85 79 89 83
rect 93 79 97 83
rect 101 79 105 83
rect 109 79 113 83
rect 117 79 121 83
rect 125 79 129 83
rect 133 79 137 83
<< nsubstratencontact >>
rect 29 1 33 5
rect 37 1 41 5
rect 45 1 49 5
rect 53 1 57 5
rect 61 1 65 5
rect 69 1 73 5
rect 77 1 81 5
rect 85 1 89 5
rect 93 1 97 5
rect 101 1 105 5
rect 109 1 113 5
rect 117 1 121 5
rect 125 1 129 5
rect 133 1 137 5
<< polysilicon >>
rect 33 75 35 77
rect 38 75 40 77
rect 54 75 56 77
rect 59 75 61 77
rect 67 75 69 77
rect 72 75 74 77
rect 81 75 83 77
rect 97 75 99 77
rect 102 75 104 77
rect 110 75 112 77
rect 115 75 117 77
rect 124 75 126 77
rect 129 75 131 77
rect 33 64 35 65
rect 38 64 40 65
rect 54 64 56 65
rect 33 62 40 64
rect 44 62 56 64
rect 33 58 35 62
rect 33 32 35 54
rect 44 46 46 62
rect 59 58 61 65
rect 54 56 61 58
rect 67 51 69 65
rect 72 62 74 65
rect 72 58 73 62
rect 72 54 74 58
rect 72 52 78 54
rect 58 49 69 51
rect 44 42 48 46
rect 44 32 46 42
rect 58 40 60 49
rect 68 41 69 45
rect 76 42 78 52
rect 60 36 61 37
rect 58 35 61 36
rect 33 30 40 32
rect 44 30 56 32
rect 33 29 35 30
rect 38 29 40 30
rect 54 29 56 30
rect 59 29 61 35
rect 67 29 69 41
rect 72 40 78 42
rect 72 29 74 40
rect 81 36 83 65
rect 97 64 99 65
rect 87 62 99 64
rect 87 46 89 62
rect 102 58 104 65
rect 97 56 104 58
rect 110 51 112 65
rect 101 49 112 51
rect 115 62 117 65
rect 124 64 126 65
rect 129 64 131 65
rect 124 62 131 64
rect 115 58 116 62
rect 101 46 103 49
rect 82 32 83 36
rect 81 29 83 32
rect 89 32 91 42
rect 101 37 103 42
rect 111 41 112 45
rect 101 35 104 37
rect 89 30 99 32
rect 97 29 99 30
rect 102 29 104 35
rect 110 29 112 41
rect 115 29 117 58
rect 124 36 126 62
rect 125 32 126 36
rect 124 30 131 32
rect 124 29 126 30
rect 129 29 131 30
rect 33 7 35 9
rect 38 7 40 9
rect 54 7 56 9
rect 59 7 61 9
rect 67 7 69 9
rect 72 7 74 9
rect 81 7 83 9
rect 97 7 99 9
rect 102 7 104 9
rect 110 7 112 9
rect 115 7 117 9
rect 124 7 126 9
rect 129 7 131 9
<< polycontact >>
rect 33 54 37 58
rect 50 54 54 58
rect 73 58 77 62
rect 48 42 52 46
rect 64 41 68 45
rect 56 36 60 40
rect 93 54 97 58
rect 116 58 120 62
rect 87 42 91 46
rect 99 42 103 46
rect 78 32 82 36
rect 107 41 111 45
rect 121 32 125 36
<< metal1 >>
rect 18 83 139 84
rect 18 79 29 83
rect 33 79 37 83
rect 41 79 45 83
rect 49 79 53 83
rect 57 79 61 83
rect 65 79 69 83
rect 73 79 77 83
rect 81 79 85 83
rect 89 79 93 83
rect 97 79 101 83
rect 105 79 109 83
rect 113 79 117 83
rect 121 79 125 83
rect 129 79 133 83
rect 137 79 139 83
rect 18 78 139 79
rect 28 75 32 78
rect 49 75 53 78
rect 75 75 80 78
rect 92 75 96 78
rect 118 75 123 78
rect 22 54 33 58
rect 22 32 25 54
rect 41 36 45 65
rect 63 55 66 65
rect 84 62 88 65
rect 77 58 88 62
rect 63 52 82 55
rect 78 36 82 52
rect 41 32 56 36
rect 63 32 78 36
rect 85 46 88 58
rect 106 55 109 65
rect 132 62 136 65
rect 120 58 136 62
rect 106 52 125 55
rect 85 42 87 46
rect 41 29 45 32
rect 63 29 66 32
rect 85 29 88 42
rect 121 36 125 52
rect 106 32 121 36
rect 106 29 109 32
rect 132 29 136 58
rect 28 6 32 9
rect 49 6 53 9
rect 75 6 80 9
rect 92 6 96 9
rect 118 6 123 9
rect 18 5 139 6
rect 18 1 29 5
rect 33 1 37 5
rect 41 1 45 5
rect 49 1 53 5
rect 57 1 61 5
rect 65 1 69 5
rect 73 1 77 5
rect 81 1 85 5
rect 89 1 93 5
rect 97 1 101 5
rect 105 1 109 5
rect 113 1 117 5
rect 121 1 125 5
rect 129 1 133 5
rect 137 1 139 5
rect 18 0 139 1
<< m2contact >>
rect 33 58 37 62
rect 50 58 54 62
rect 48 46 52 50
rect 64 45 68 49
rect 56 32 60 36
rect 93 50 97 54
rect 95 42 99 46
rect 107 45 111 49
<< metal2 >>
rect 22 71 30 75
rect 26 50 30 71
rect 37 58 50 62
rect 54 58 60 62
rect 26 46 48 50
rect 56 49 60 58
rect 97 50 111 54
rect 107 49 111 50
rect 56 45 64 49
rect 68 46 88 49
rect 68 45 95 46
rect 84 42 95 45
rect 107 36 111 45
rect 60 32 111 36
<< labels >>
rlabel metal2 24 73 24 73 1 D
rlabel metal1 23 45 23 45 3 clk_b
rlabel metal1 43 45 43 45 1 clk
rlabel metal1 135 45 135 45 7 Q
<< end >>
