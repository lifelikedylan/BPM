magic
tech scmos
timestamp 1542725905
<< metal1 >>
rect -8 -2 -7 2
rect -3 -2 3 2
rect 7 -2 8 2
<< m2contact >>
rect -7 -2 -3 2
rect 3 -2 7 2
<< metal2 >>
rect -8 -2 -7 2
rect -3 -2 3 2
rect 7 -2 8 2
<< end >>
