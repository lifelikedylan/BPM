magic
tech scmos
magscale 1 2
timestamp 1542729052
<< metal1 >>
rect 2044 7812 7956 7908
rect 1996 7686 2140 7796
rect 2164 7692 7836 7788
rect 7860 7686 8004 7796
rect 1996 7674 8004 7686
rect 1996 7604 2140 7674
rect 7860 7604 8004 7674
rect 2164 7474 7836 7486
rect 4453 7407 5531 7413
rect 2044 7274 7956 7286
rect 1996 7086 2260 7196
rect 7740 7086 8004 7196
rect 1996 7074 8004 7086
rect 1996 7004 2260 7074
rect 4549 7007 4651 7013
rect 4645 6993 4651 7007
rect 7740 7004 8004 7074
rect 4408 6987 4619 6993
rect 4645 6987 4824 6993
rect 4613 6973 4619 6987
rect 4392 6967 4411 6973
rect 4613 6967 4840 6973
rect 4325 6947 4376 6953
rect 4856 6947 5035 6953
rect 5125 6947 5256 6953
rect 5029 6933 5035 6947
rect 5029 6927 5240 6933
rect 2044 6874 7956 6886
rect 4597 6827 4824 6833
rect 4597 6813 4603 6827
rect 4229 6807 4344 6813
rect 4392 6807 4603 6813
rect 4840 6807 5035 6813
rect 5157 6807 5192 6813
rect 5240 6810 5560 6813
rect 5240 6807 5563 6810
rect 5656 6807 5707 6813
rect 5029 6793 5035 6807
rect 5029 6787 5208 6793
rect 5557 6787 5563 6807
rect 5608 6787 5627 6793
rect 5701 6787 5707 6807
rect 4392 6767 4411 6773
rect 2164 6674 7836 6686
rect 5077 6587 5208 6593
rect 5557 6587 5672 6593
rect 5781 6587 5896 6593
rect 6277 6587 6296 6593
rect 5781 6573 5787 6587
rect 4181 6567 4360 6573
rect 4773 6567 4811 6573
rect 4853 6567 5224 6573
rect 5688 6567 5787 6573
rect 5928 6567 6011 6573
rect 6165 6567 6312 6573
rect 4181 6553 4187 6567
rect 3861 6547 4187 6553
rect 4392 6547 4795 6553
rect 4805 6550 4811 6567
rect 6165 6553 6171 6567
rect 5240 6547 5451 6553
rect 5765 6547 5896 6553
rect 5944 6547 6171 6553
rect 6328 6547 6731 6553
rect 2044 6474 7956 6486
rect 4440 6427 4459 6433
rect 4792 6427 4811 6433
rect 3429 6407 3832 6413
rect 3925 6407 4424 6413
rect 4853 6407 5128 6413
rect 5397 6407 5432 6413
rect 5480 6407 5691 6413
rect 5701 6407 5928 6413
rect 3848 6387 3867 6393
rect 4437 6387 4760 6393
rect 5144 6387 5227 6393
rect 5429 6387 5448 6393
rect 5685 6373 5691 6407
rect 5685 6367 5928 6373
rect 2164 6274 7836 6286
rect 3480 6187 3531 6193
rect 4168 6167 4187 6173
rect 4581 6167 4744 6173
rect 5589 6167 5624 6173
rect 5672 6167 5883 6173
rect 3480 6147 3819 6153
rect 3845 6147 4152 6153
rect 4709 6147 4728 6153
rect 4952 6147 5160 6153
rect 5384 6147 5611 6153
rect 5877 6147 5883 6167
rect 6005 6147 6232 6153
rect 4053 6127 4136 6133
rect 5672 6127 5947 6133
rect 5973 6127 6216 6133
rect 2044 6074 7956 6086
rect 3509 6007 3992 6013
rect 4040 6007 4059 6013
rect 4453 6007 4504 6013
rect 4709 6007 4936 6013
rect 5173 6007 5352 6013
rect 4024 5987 4187 5993
rect 4520 5987 4891 5993
rect 4952 5987 4971 5993
rect 5317 5987 5336 5993
rect 5365 5987 5371 6030
rect 5381 6007 5672 6013
rect 5768 6007 5931 6013
rect 5720 5987 5739 5993
rect 3909 5967 3992 5973
rect 4536 5967 4555 5973
rect 4549 5947 4555 5967
rect 5925 5953 5931 6007
rect 5941 5967 5959 5973
rect 6008 5967 6027 5973
rect 5925 5947 5992 5953
rect 2164 5874 7836 5886
rect 3909 5787 4235 5793
rect 5912 5787 6027 5793
rect 4229 5773 4235 5787
rect 4229 5767 4424 5773
rect 4472 5767 4587 5773
rect 5061 5754 5067 5773
rect 3461 5747 3512 5753
rect 3845 5747 4440 5753
rect 4792 5747 4971 5753
rect 5189 5747 5384 5753
rect 5608 5747 5803 5753
rect 5829 5747 5864 5753
rect 5912 5747 6075 5753
rect 6216 5747 6363 5753
rect 6488 5747 6571 5753
rect 4661 5727 4776 5733
rect 5829 5713 5835 5747
rect 6069 5733 6075 5747
rect 6357 5733 6363 5747
rect 6069 5727 6200 5733
rect 6357 5727 6472 5733
rect 5621 5707 5835 5713
rect 2044 5674 7956 5686
rect 6021 5647 6155 5653
rect 6149 5633 6155 5647
rect 4936 5627 5051 5633
rect 5365 5627 5419 5633
rect 5976 5627 6107 5633
rect 6149 5627 6184 5633
rect 6552 5627 6571 5633
rect 3896 5607 4203 5613
rect 4472 5607 4555 5613
rect 5077 5607 5192 5613
rect 5365 5593 5371 5627
rect 6101 5613 6107 5627
rect 3461 5587 3864 5593
rect 4213 5587 4424 5593
rect 4488 5587 4523 5593
rect 5208 5587 5371 5593
rect 5397 5593 5403 5613
rect 5877 5593 5883 5613
rect 5960 5607 5995 5613
rect 6101 5607 6200 5613
rect 6469 5607 6520 5613
rect 5397 5587 5544 5593
rect 5877 5587 5940 5593
rect 6552 5587 6603 5593
rect 3896 5567 3915 5573
rect 5224 5567 5259 5573
rect 5509 5567 5528 5573
rect 2164 5474 7836 5486
rect 4549 5367 4760 5373
rect 5080 5367 5147 5373
rect 4053 5347 4232 5353
rect 4405 5347 4520 5353
rect 4776 5347 5032 5353
rect 5157 5347 5515 5353
rect 5528 5347 5755 5353
rect 5768 5347 5867 5353
rect 5893 5347 6280 5353
rect 6376 5347 6776 5353
rect 5893 5333 5899 5347
rect 4485 5327 4504 5333
rect 5253 5327 5288 5333
rect 5493 5327 5511 5333
rect 5717 5327 5752 5333
rect 5781 5327 5899 5333
rect 2044 5274 7956 5286
rect 6520 5227 6571 5233
rect 4408 5207 4491 5213
rect 4744 5207 4763 5213
rect 4965 5207 5000 5213
rect 5352 5207 5499 5213
rect 5861 5207 5928 5213
rect 6504 5207 6827 5213
rect 4661 5187 4712 5193
rect 6437 5187 6472 5193
rect 4744 5167 4763 5173
rect 4757 5086 4763 5167
rect 2164 5074 7836 5086
rect 4619 5025 6571 5037
rect 4643 5001 6547 5013
rect 5676 4987 5739 4993
rect 6145 4987 6187 4993
rect 3816 4967 3851 4973
rect 4117 4967 4152 4973
rect 4677 4967 4891 4973
rect 5013 4967 5046 4973
rect 5205 4967 5234 4973
rect 4677 4953 4683 4967
rect 4184 4947 4459 4953
rect 4520 4947 4683 4953
rect 4800 4950 4806 4967
rect 5040 4950 5046 4967
rect 5228 4950 5234 4967
rect 5249 4967 5323 4973
rect 5489 4967 5659 4973
rect 5249 4950 5255 4967
rect 5489 4950 5495 4967
rect 5676 4950 5682 4987
rect 5697 4967 5755 4973
rect 5893 4967 5942 4973
rect 5697 4950 5703 4967
rect 5936 4950 5942 4967
rect 6145 4950 6151 4987
rect 6181 4983 6187 4987
rect 6357 4987 6875 4993
rect 6357 4983 6363 4987
rect 6181 4977 6363 4983
rect 6385 4967 6603 4973
rect 6385 4950 6391 4967
rect 2044 4874 4631 4886
rect 6559 4874 7956 4886
rect 4437 4707 4667 4713
rect 4661 4693 4667 4707
rect 4800 4693 4806 4700
rect 5040 4693 5046 4700
rect 5248 4693 5254 4700
rect 4661 4687 4806 4693
rect 4837 4687 4875 4693
rect 2164 4674 4655 4686
rect 4869 4683 4875 4687
rect 5013 4687 5046 4693
rect 5221 4687 5254 4693
rect 5013 4683 5019 4687
rect 4869 4677 5019 4683
rect 5285 4677 5467 4683
rect 5285 4673 5291 4677
rect 5141 4667 5291 4673
rect 5461 4673 5467 4677
rect 5488 4673 5494 4700
rect 5696 4673 5702 4700
rect 5937 4693 5943 4700
rect 6144 4693 6150 4700
rect 5937 4687 5995 4693
rect 6117 4687 6150 4693
rect 5461 4667 5494 4673
rect 5525 4667 5702 4673
rect 6385 4673 6391 4700
rect 6405 4693 6411 4705
rect 6405 4687 6523 4693
rect 6535 4674 7836 4686
rect 6385 4667 6411 4673
rect 4643 4643 6547 4655
rect 4619 4619 6571 4631
rect 4104 4607 4123 4613
rect 3797 4587 3816 4593
rect 2044 4474 7956 4486
rect 6872 4407 7675 4413
rect 6549 4387 6840 4393
rect 4293 4367 4312 4373
rect 6549 4353 6555 4387
rect 6328 4347 6555 4353
rect 2164 4274 7836 4286
rect 5720 4207 5947 4213
rect 5413 4187 5432 4193
rect 5941 4173 5947 4207
rect 5941 4167 6088 4173
rect 6120 4147 6283 4153
rect 2044 4074 7956 4086
rect 5061 3967 5080 3973
rect 5829 3967 5848 3973
rect 5368 3947 5387 3953
rect 6136 3947 6171 3953
rect 2164 3874 7836 3886
rect 5381 3767 5400 3773
rect 5765 3753 5771 3773
rect 6632 3767 7115 3773
rect 5432 3747 5771 3753
rect 2044 3674 7956 3686
rect 5845 3607 5960 3613
rect 5992 3587 6171 3593
rect 2164 3474 7836 3486
rect 2044 3274 7956 3286
rect 6293 3167 7979 3173
rect 2164 3074 7836 3086
rect 6597 2927 7307 2933
rect 2044 2874 7956 2886
rect 2164 2674 7836 2686
rect 2044 2474 7956 2486
rect 5941 2307 7851 2313
rect 2164 2274 7836 2286
rect 2164 2172 7836 2268
rect 2044 2052 7956 2148
rect 7685 2027 7883 2033
<< metal2 >>
rect 2044 2052 2140 7908
rect 2164 2172 2260 7788
rect 4357 6987 4411 6993
rect 4213 6807 4235 6813
rect 4325 6807 4331 6953
rect 4133 6727 4155 6733
rect 3813 6427 3835 6433
rect 3429 6113 3435 6413
rect 3861 6387 3867 6553
rect 3957 6507 3963 6533
rect 3925 6407 3931 6433
rect 3445 6167 3499 6173
rect 3429 6107 3451 6113
rect 3445 5793 3451 6107
rect 3493 6013 3499 6167
rect 3525 6153 3531 6193
rect 3525 6147 3547 6153
rect 3813 6147 3835 6153
rect 3493 6007 3515 6013
rect 3445 5787 3467 5793
rect 3461 5587 3467 5787
rect 3493 5733 3499 6007
rect 3541 5833 3547 6147
rect 3525 5827 3547 5833
rect 3525 5767 3531 5827
rect 3541 5733 3547 5793
rect 3493 5727 3547 5733
rect 3045 4327 3051 5573
rect 3525 3727 3531 5213
rect 3797 4947 3803 6133
rect 3845 5607 3851 6153
rect 3909 5567 3915 5973
rect 4053 5347 4059 6133
rect 4101 5567 4107 6513
rect 3797 4587 3803 4683
rect 3845 4407 3851 4973
rect 4117 4933 4123 4973
rect 4101 4927 4123 4933
rect 4101 4653 4107 4927
rect 4101 4647 4123 4653
rect 3909 4527 3915 4553
rect 3941 4527 3947 4633
rect 4117 4607 4123 4647
rect 4149 4287 4155 6727
rect 4213 6433 4219 6807
rect 4357 6787 4363 6987
rect 4389 6587 4395 6813
rect 4405 6767 4411 6973
rect 4341 6567 4395 6573
rect 4213 6427 4235 6433
rect 4181 5987 4187 6413
rect 4229 5973 4235 6427
rect 4341 6107 4347 6553
rect 4389 6393 4395 6567
rect 4389 6387 4443 6393
rect 4213 5967 4235 5973
rect 4213 5747 4219 5967
rect 4453 5933 4459 7413
rect 4549 6193 4555 7013
rect 4773 6567 4779 6833
rect 4789 6587 4859 6593
rect 4789 6547 4795 6587
rect 4821 6567 4859 6573
rect 4773 6373 4779 6413
rect 4533 6187 4555 6193
rect 4757 6367 4779 6373
rect 4533 5993 4539 6187
rect 4581 6013 4587 6173
rect 4757 6167 4763 6367
rect 4805 6207 4811 6433
rect 4853 6407 4859 6553
rect 4917 6207 4923 8000
rect 5525 7407 5531 8000
rect 5125 6833 5131 6953
rect 6117 6947 6123 8000
rect 5221 6927 5243 6933
rect 5109 6827 5131 6833
rect 5109 6633 5115 6827
rect 5109 6627 5131 6633
rect 5077 6487 5083 6593
rect 4581 6007 4603 6013
rect 4709 6007 4715 6153
rect 4533 5987 4555 5993
rect 4453 5927 4507 5933
rect 4437 5793 4443 5833
rect 4429 5787 4443 5793
rect 4405 5733 4411 5773
rect 4197 5607 4203 5733
rect 4389 5727 4411 5733
rect 4389 5593 4395 5727
rect 4429 5653 4435 5787
rect 4501 5773 4507 5927
rect 4501 5767 4523 5773
rect 4453 5727 4475 5733
rect 4429 5647 4443 5653
rect 4437 5607 4443 5647
rect 4213 5453 4219 5593
rect 4389 5587 4411 5593
rect 4453 5587 4459 5727
rect 4181 5447 4219 5453
rect 4213 5327 4219 5447
rect 4405 5347 4411 5587
rect 4469 5333 4475 5613
rect 4517 5527 4523 5767
rect 4549 5607 4555 5987
rect 4597 5813 4603 6007
rect 4581 5807 4603 5813
rect 4581 5767 4587 5807
rect 4533 5367 4539 5393
rect 4549 5333 4555 5373
rect 4661 5353 4667 5733
rect 4389 5327 4475 5333
rect 4485 5327 4555 5333
rect 4645 5347 4667 5353
rect 4389 4907 4395 5327
rect 4485 5207 4491 5327
rect 4645 5233 4651 5347
rect 4741 5333 4747 6113
rect 4805 5767 4811 6173
rect 4933 6107 4939 6133
rect 4885 5967 4891 5993
rect 4917 5607 4923 6033
rect 4965 5967 4971 5993
rect 5061 5767 5067 6413
rect 5125 6393 5131 6627
rect 5157 6567 5163 6813
rect 5237 6573 5243 6773
rect 5557 6587 5563 6793
rect 5221 6567 5243 6573
rect 5429 6567 5467 6573
rect 5109 6387 5131 6393
rect 5221 6387 5227 6567
rect 5109 6053 5115 6387
rect 5397 6373 5403 6413
rect 5157 6193 5163 6373
rect 5381 6367 5403 6373
rect 5381 6233 5387 6367
rect 5381 6227 5403 6233
rect 5141 6187 5163 6193
rect 5141 6093 5147 6187
rect 5141 6087 5155 6093
rect 5109 6047 5131 6053
rect 5125 6007 5131 6047
rect 5149 5993 5155 6087
rect 5173 6007 5179 6173
rect 5189 6147 5195 6173
rect 5149 5987 5163 5993
rect 5109 5767 5115 5793
rect 4965 5627 4971 5753
rect 4693 5327 4795 5333
rect 4645 5227 4667 5233
rect 4661 5187 4667 5227
rect 4693 5207 4699 5327
rect 4453 4947 4459 4993
rect 4405 4707 4443 4713
rect 4341 4387 4347 4413
rect 4405 4407 4411 4707
rect 4485 4687 4491 4973
rect 4293 4277 4299 4373
rect 4437 4287 4443 4433
rect 4597 4347 4603 4693
rect 4619 4619 4631 5037
rect 4643 4643 4655 5013
rect 4699 4947 4719 5037
rect 4757 4953 4763 5213
rect 4757 4947 4786 4953
rect 4821 4947 4827 5033
rect 4885 4967 4891 5493
rect 5045 5353 5051 5633
rect 5077 5567 5083 5613
rect 5157 5433 5163 5987
rect 5253 5793 5259 6173
rect 5365 6073 5371 6133
rect 5365 6067 5387 6073
rect 5317 5987 5323 6013
rect 5381 6007 5387 6067
rect 5397 5993 5403 6227
rect 5429 6067 5435 6567
rect 5445 6533 5451 6553
rect 5461 6547 5467 6567
rect 5445 6527 5483 6533
rect 5477 6513 5483 6527
rect 5477 6507 5499 6513
rect 5621 6407 5627 6793
rect 5701 6407 5707 6793
rect 5477 6253 5483 6373
rect 5477 6247 5499 6253
rect 5477 6107 5483 6247
rect 5589 6007 5595 6173
rect 5605 6133 5611 6153
rect 5637 6147 5643 6173
rect 5605 6127 5675 6133
rect 5765 6007 5771 6553
rect 5957 6387 5963 6553
rect 6005 6433 6011 6573
rect 6005 6427 6027 6433
rect 5365 5987 5403 5993
rect 5365 5793 5371 5987
rect 5189 5727 5195 5753
rect 5221 5593 5227 5793
rect 5253 5787 5275 5793
rect 5269 5613 5275 5787
rect 5141 5427 5163 5433
rect 5205 5587 5227 5593
rect 5253 5607 5275 5613
rect 5349 5787 5371 5793
rect 5141 5367 5147 5427
rect 4965 5207 4971 5353
rect 5045 5347 5099 5353
rect 5157 5347 5163 5393
rect 5093 5207 5099 5347
rect 5045 5013 5051 5193
rect 4907 4955 4939 5013
rect 5045 5007 5067 5013
rect 5013 4967 5019 4993
rect 5061 4947 5067 5007
rect 5127 4954 5167 5037
rect 5205 4967 5211 5587
rect 5253 5327 5259 5607
rect 5349 5593 5355 5787
rect 5397 5607 5403 5773
rect 5413 5627 5419 5773
rect 5589 5713 5595 5733
rect 5589 5707 5627 5713
rect 5717 5673 5723 5713
rect 5685 5667 5723 5673
rect 5349 5587 5371 5593
rect 5365 5413 5371 5587
rect 5509 5527 5515 5573
rect 5365 5407 5387 5413
rect 5333 5227 5339 5393
rect 5381 5253 5387 5407
rect 5541 5353 5547 5373
rect 5509 5347 5547 5353
rect 5365 5247 5387 5253
rect 5365 5207 5371 5247
rect 5493 5207 5499 5333
rect 5557 5147 5563 5613
rect 5685 5373 5691 5667
rect 5685 5367 5723 5373
rect 5717 5327 5723 5367
rect 5317 4867 5323 4973
rect 5355 4954 5387 5013
rect 5509 4947 5515 5013
rect 5575 4954 5615 5037
rect 5733 4987 5739 5993
rect 5797 5727 5803 5753
rect 5877 5607 5883 6153
rect 5941 5967 5947 6133
rect 5973 6127 5979 6413
rect 6021 6193 6027 6427
rect 6005 6187 6027 6193
rect 6005 6147 6011 6187
rect 5973 5987 5979 6033
rect 6021 5647 6027 5973
rect 5989 5553 5995 5613
rect 5989 5547 6027 5553
rect 5749 5347 5787 5353
rect 5781 5327 5787 5347
rect 5861 5207 5867 5353
rect 6021 5207 6027 5547
rect 5973 5033 5979 5193
rect 5957 5027 5979 5033
rect 5653 4933 5659 4973
rect 5749 4947 5755 4973
rect 5803 4954 5835 5013
rect 5653 4927 5771 4933
rect 5893 4927 5899 4973
rect 5957 4947 5963 5027
rect 6023 4954 6063 5037
rect 6149 4953 6155 5393
rect 6261 5327 6267 5353
rect 6277 5147 6283 6593
rect 6325 6527 6331 6553
rect 6725 6547 6731 8000
rect 6389 6407 6411 6413
rect 6325 5367 6331 5393
rect 6405 5213 6411 6407
rect 6453 5673 6459 5733
rect 6453 5667 6475 5673
rect 6469 5607 6475 5667
rect 6501 5587 6507 5773
rect 6565 5593 6571 5753
rect 6549 5587 6571 5593
rect 6549 5333 6555 5587
rect 6597 5347 6603 5593
rect 6549 5327 6571 5333
rect 6789 5327 6795 5373
rect 6565 5227 6571 5327
rect 6389 5207 6411 5213
rect 6821 5207 6827 5373
rect 6389 5073 6395 5207
rect 6389 5067 6411 5073
rect 6405 5027 6411 5067
rect 6251 4954 6283 5013
rect 6437 4973 6443 5193
rect 6405 4967 6443 4973
rect 6263 4953 6271 4954
rect 6124 4947 6155 4953
rect 6405 4947 6411 4967
rect 6471 4947 6491 5037
rect 5397 4867 5419 4873
rect 5413 4833 5419 4867
rect 5397 4827 5419 4833
rect 4699 4619 4719 4713
rect 4837 4527 4843 4693
rect 4919 4643 4927 4707
rect 5397 4693 5403 4827
rect 5765 4807 5771 4927
rect 5813 4693 5819 4813
rect 5093 4407 5115 4413
rect 5109 4153 5115 4407
rect 5125 4277 5131 4373
rect 5093 4147 5115 4153
rect 5093 4033 5099 4147
rect 5141 4113 5147 4673
rect 5221 4407 5227 4693
rect 5397 4687 5419 4693
rect 5157 4307 5163 4393
rect 5173 4127 5179 4293
rect 5253 4287 5259 4433
rect 5413 4307 5419 4687
rect 5765 4687 5819 4693
rect 5413 4187 5419 4283
rect 5461 4167 5467 4193
rect 5525 4147 5531 4673
rect 5141 4107 5179 4113
rect 5093 4027 5115 4033
rect 5109 3987 5115 4027
rect 5173 4007 5179 4107
rect 5205 4027 5211 4133
rect 5525 4087 5531 4133
rect 5557 4087 5563 4129
rect 5061 3877 5067 3973
rect 5381 3767 5387 3953
rect 5765 3707 5771 4687
rect 5845 4213 5851 4873
rect 6277 4733 6283 4873
rect 6277 4727 6299 4733
rect 5829 4207 5851 4213
rect 5829 4013 5835 4207
rect 5829 4007 5851 4013
rect 5845 3973 5851 4007
rect 5829 3877 5835 3973
rect 5845 3967 5859 3973
rect 5877 3967 5883 4193
rect 5941 4007 5947 4053
rect 5973 4027 5979 4133
rect 5989 4067 5995 4693
rect 6117 4673 6123 4693
rect 6117 4667 6139 4673
rect 6133 4407 6139 4667
rect 6263 4643 6271 4707
rect 6293 4633 6299 4727
rect 6277 4627 6299 4633
rect 6037 4277 6043 4373
rect 6069 3967 6075 4393
rect 6165 4127 6171 4433
rect 6277 4153 6283 4627
rect 6277 4147 6299 4153
rect 5853 3873 5859 3967
rect 5845 3867 5859 3873
rect 5845 3607 5851 3867
rect 5941 2307 5947 3613
rect 6165 3587 6171 3953
rect 6293 3167 6299 4147
rect 6405 4027 6411 4673
rect 6471 4619 6491 4713
rect 6517 2147 6523 4693
rect 6535 4643 6547 5013
rect 6559 4619 6571 5037
rect 6597 4933 6603 4973
rect 6597 4927 6619 4933
rect 6613 4613 6619 4927
rect 6597 4607 6619 4613
rect 6597 2927 6603 4607
rect 6869 4407 6875 4993
rect 7669 4407 7691 4413
rect 6917 4007 6923 4033
rect 6949 4027 6955 4133
rect 6821 3877 6827 3973
rect 6853 3967 6859 3993
rect 7109 3767 7115 3953
rect 6677 2147 6707 2153
rect 6701 2000 6707 2147
rect 7301 2000 7307 2933
rect 7685 2027 7691 4407
rect 7740 2172 7836 7788
rect 7845 2307 7851 2513
rect 7860 2052 7956 7908
rect 7973 3107 7979 3173
rect 7877 2027 7907 2033
rect 7901 2000 7907 2027
<< metal3 >>
rect 4526 9530 4880 9948
rect 5110 9558 5464 9976
rect 5732 9558 6086 9976
rect 6308 9548 6662 9966
rect 104 7452 458 7870
rect 9544 7498 9898 7916
rect 66 6924 420 7342
rect 6115 6935 6125 6955
rect 5235 6925 6125 6935
rect 9572 6878 9926 7296
rect 1993 6725 4141 6735
rect 94 6302 448 6720
rect 5539 6525 6333 6535
rect 5539 6515 5549 6525
rect 3955 6505 4493 6515
rect 5491 6505 5549 6515
rect 4483 6495 4493 6505
rect 4483 6485 5085 6495
rect 3827 6425 3933 6435
rect 5619 6405 6397 6415
rect 5491 6245 5981 6255
rect 4803 6165 4813 6215
rect 4915 6205 5197 6215
rect 5187 6175 5197 6205
rect 5187 6165 5261 6175
rect 5635 6165 5773 6175
rect 3827 6145 5197 6155
rect 84 5708 438 6126
rect 1993 6125 3805 6135
rect 5299 6125 5437 6135
rect 5299 6115 5309 6125
rect 4339 6105 4397 6115
rect 4387 6095 4397 6105
rect 4691 6105 4909 6115
rect 4931 6105 5309 6115
rect 5427 6115 5437 6125
rect 5427 6105 5485 6115
rect 4691 6095 4701 6105
rect 4387 6085 4701 6095
rect 4899 6075 4909 6105
rect 4899 6065 5437 6075
rect 5587 6025 5981 6035
rect 4803 6005 5325 6015
rect 4883 5965 4973 5975
rect 5075 5845 5213 5855
rect 5075 5835 5085 5845
rect 4435 5825 5085 5835
rect 5203 5835 5213 5845
rect 5203 5825 5261 5835
rect 5107 5785 5229 5795
rect 4195 5725 5197 5735
rect 5795 5725 6509 5735
rect 4051 5685 4173 5695
rect 4163 5675 4173 5685
rect 4611 5685 4669 5695
rect 4611 5675 4621 5685
rect 4163 5665 4621 5675
rect 4803 5585 5037 5595
rect 4803 5575 4813 5585
rect 3043 5565 4813 5575
rect 5027 5575 5037 5585
rect 5027 5565 5085 5575
rect 1993 5525 2157 5535
rect 4515 5525 4573 5535
rect 76 5096 430 5514
rect 2147 5455 2157 5525
rect 4563 5515 4573 5525
rect 4835 5525 5517 5535
rect 4835 5515 4845 5525
rect 4563 5505 4845 5515
rect 5507 5505 8007 5515
rect 4883 5485 4941 5495
rect 4931 5475 4941 5485
rect 5507 5475 5517 5505
rect 4931 5465 5517 5475
rect 2147 5445 4189 5455
rect 4531 5385 5165 5395
rect 5331 5385 5565 5395
rect 6147 5385 6333 5395
rect 6259 5325 6797 5335
rect 5251 5245 5341 5255
rect 5251 5235 5261 5245
rect 3523 5225 5261 5235
rect 3523 5205 3533 5225
rect 5555 5145 6285 5155
rect 9580 5096 9934 5514
rect 5667 5025 6093 5035
rect 5667 5015 5677 5025
rect 5507 5005 5677 5015
rect 6083 5015 6093 5025
rect 6403 5015 6413 5035
rect 6083 5005 6413 5015
rect 4451 4985 5517 4995
rect 5507 4955 5517 4985
rect 5731 4985 6029 4995
rect 5731 4975 5741 4985
rect 5699 4965 5741 4975
rect 6019 4975 6029 4985
rect 6019 4965 6061 4975
rect 5699 4955 5709 4965
rect 5507 4945 5709 4955
rect 5747 4945 5933 4955
rect 84 4522 438 4940
rect 1993 4925 2125 4935
rect 2115 4915 2125 4925
rect 2115 4905 4397 4915
rect 5891 4875 5901 4935
rect 5315 4865 5405 4875
rect 5843 4865 5901 4875
rect 5923 4855 5933 4945
rect 6051 4915 6061 4965
rect 6051 4905 8007 4915
rect 6227 4865 6285 4875
rect 6227 4855 6237 4865
rect 5923 4845 6237 4855
rect 5763 4805 5821 4815
rect 4483 4685 4605 4695
rect 3939 4625 4157 4635
rect 3907 4525 4845 4535
rect 9580 4504 9934 4922
rect 3843 4405 5101 4415
rect 1993 4325 3053 4335
rect 84 3900 438 4318
rect 5107 4305 5165 4315
rect 5411 4305 8007 4315
rect 4147 4285 5261 4295
rect 5107 4185 5885 4195
rect 5171 4125 6957 4135
rect 5523 4085 5565 4095
rect 5987 4055 5997 4075
rect 5939 4045 5997 4055
rect 6403 4025 6925 4035
rect 5875 3965 6861 3975
rect 9590 3892 9944 4310
rect 48 3316 402 3734
rect 1993 3725 3533 3735
rect 5763 3705 8007 3715
rect 9590 3298 9944 3716
rect 7971 3105 8007 3115
rect 9562 2722 9916 3140
rect 7843 2505 8007 2515
rect 6515 2145 6685 2155
rect 9552 2092 9906 2510
rect 6308 70 6662 488
rect 6892 62 7246 480
rect 7494 62 7848 480
use PADFC  PADFC_1
timestamp 949001400
transform 1 0 0 0 1 8000
box 654 -6 2006 1346
use PADNC  PADNC_0
timestamp 1084294400
transform 1 0 2000 0 1 8000
box -6 -6 606 2000
use PADNC  PADNC_1
timestamp 1084294400
transform 1 0 2600 0 1 8000
box -6 -6 606 2000
use PADNC  PADNC_2
timestamp 1084294400
transform 1 0 3200 0 1 8000
box -6 -6 606 2000
use PADNC  PADNC_3
timestamp 1084294400
transform 1 0 3800 0 1 8000
box -6 -6 606 2000
use PADINC  PADINC_0
timestamp 1084294328
transform 1 0 4400 0 1 8000
box -12 -6 606 2000
use PADINC  PADINC_1
timestamp 1084294328
transform 1 0 5000 0 1 8000
box -12 -6 606 2000
use PADINC  PADINC_2
timestamp 1084294328
transform 1 0 5600 0 1 8000
box -12 -6 606 2000
use PADINC  PADINC_3
timestamp 1084294328
transform 1 0 6200 0 1 8000
box -12 -6 606 2000
use PADNC  PADNC_4
timestamp 1084294400
transform 1 0 6800 0 1 8000
box -6 -6 606 2000
use PADNC  PADNC_5
timestamp 1084294400
transform 1 0 7400 0 1 8000
box -6 -6 606 2000
use PADFC  PADFC_0
timestamp 949001400
transform 0 1 8000 -1 0 10000
box 654 -6 2006 1346
use mult_pad_VIA0  mult_pad_VIA0_0
timestamp 1542725905
transform 1 0 2092 0 1 7860
box -48 -48 48 48
use mult_pad_VIA0  mult_pad_VIA0_1
timestamp 1542725905
transform 1 0 7908 0 1 7860
box -48 -48 48 48
use mult_pad_VIA6  mult_pad_VIA6_0
timestamp 1542725905
transform 1 0 2092 0 1 7700
box -48 -96 48 96
use mult_pad_VIA0  mult_pad_VIA0_2
timestamp 1542725905
transform 1 0 2212 0 1 7740
box -48 -48 48 48
use mult_pad_VIA0  mult_pad_VIA0_3
timestamp 1542725905
transform 1 0 7788 0 1 7740
box -48 -48 48 48
use mult_pad_VIA6  mult_pad_VIA6_1
timestamp 1542725905
transform 1 0 7908 0 1 7700
box -48 -96 48 96
use mult_pad_VIA1  mult_pad_VIA1_0
timestamp 1542725905
transform 1 0 2212 0 1 7480
box -48 -6 48 6
use PADGND  PADGND_1
timestamp 1084294269
transform 0 -1 2000 1 0 7400
box -6 -6 606 2000
use FILL  FILL_0
timestamp 1018054153
transform 1 0 2272 0 -1 7680
box -16 -6 32 210
use FILL  FILL_1
timestamp 1018054153
transform 1 0 2288 0 -1 7680
box -16 -6 32 210
use FILL  FILL_2
timestamp 1018054153
transform 1 0 2304 0 -1 7680
box -16 -6 32 210
use FILL  FILL_3
timestamp 1018054153
transform 1 0 2320 0 -1 7680
box -16 -6 32 210
use FILL  FILL_4
timestamp 1018054153
transform 1 0 2336 0 -1 7680
box -16 -6 32 210
use FILL  FILL_5
timestamp 1018054153
transform 1 0 2352 0 -1 7680
box -16 -6 32 210
use FILL  FILL_6
timestamp 1018054153
transform 1 0 2368 0 -1 7680
box -16 -6 32 210
use FILL  FILL_7
timestamp 1018054153
transform 1 0 2384 0 -1 7680
box -16 -6 32 210
use FILL  FILL_8
timestamp 1018054153
transform 1 0 2400 0 -1 7680
box -16 -6 32 210
use FILL  FILL_9
timestamp 1018054153
transform 1 0 2416 0 -1 7680
box -16 -6 32 210
use FILL  FILL_10
timestamp 1018054153
transform 1 0 2432 0 -1 7680
box -16 -6 32 210
use FILL  FILL_11
timestamp 1018054153
transform 1 0 2448 0 -1 7680
box -16 -6 32 210
use FILL  FILL_12
timestamp 1018054153
transform 1 0 2464 0 -1 7680
box -16 -6 32 210
use FILL  FILL_13
timestamp 1018054153
transform 1 0 2480 0 -1 7680
box -16 -6 32 210
use FILL  FILL_14
timestamp 1018054153
transform 1 0 2496 0 -1 7680
box -16 -6 32 210
use FILL  FILL_15
timestamp 1018054153
transform 1 0 2512 0 -1 7680
box -16 -6 32 210
use FILL  FILL_16
timestamp 1018054153
transform 1 0 2528 0 -1 7680
box -16 -6 32 210
use FILL  FILL_17
timestamp 1018054153
transform 1 0 2544 0 -1 7680
box -16 -6 32 210
use FILL  FILL_18
timestamp 1018054153
transform 1 0 2560 0 -1 7680
box -16 -6 32 210
use FILL  FILL_19
timestamp 1018054153
transform 1 0 2576 0 -1 7680
box -16 -6 32 210
use FILL  FILL_20
timestamp 1018054153
transform 1 0 2592 0 -1 7680
box -16 -6 32 210
use FILL  FILL_21
timestamp 1018054153
transform 1 0 2608 0 -1 7680
box -16 -6 32 210
use FILL  FILL_22
timestamp 1018054153
transform 1 0 2624 0 -1 7680
box -16 -6 32 210
use FILL  FILL_23
timestamp 1018054153
transform 1 0 2640 0 -1 7680
box -16 -6 32 210
use FILL  FILL_24
timestamp 1018054153
transform 1 0 2656 0 -1 7680
box -16 -6 32 210
use FILL  FILL_25
timestamp 1018054153
transform 1 0 2672 0 -1 7680
box -16 -6 32 210
use FILL  FILL_26
timestamp 1018054153
transform 1 0 2688 0 -1 7680
box -16 -6 32 210
use FILL  FILL_27
timestamp 1018054153
transform 1 0 2704 0 -1 7680
box -16 -6 32 210
use FILL  FILL_28
timestamp 1018054153
transform 1 0 2720 0 -1 7680
box -16 -6 32 210
use FILL  FILL_29
timestamp 1018054153
transform 1 0 2736 0 -1 7680
box -16 -6 32 210
use FILL  FILL_30
timestamp 1018054153
transform 1 0 2752 0 -1 7680
box -16 -6 32 210
use FILL  FILL_31
timestamp 1018054153
transform 1 0 2768 0 -1 7680
box -16 -6 32 210
use FILL  FILL_32
timestamp 1018054153
transform 1 0 2784 0 -1 7680
box -16 -6 32 210
use FILL  FILL_33
timestamp 1018054153
transform 1 0 2800 0 -1 7680
box -16 -6 32 210
use FILL  FILL_34
timestamp 1018054153
transform 1 0 2816 0 -1 7680
box -16 -6 32 210
use FILL  FILL_35
timestamp 1018054153
transform 1 0 2832 0 -1 7680
box -16 -6 32 210
use FILL  FILL_36
timestamp 1018054153
transform 1 0 2848 0 -1 7680
box -16 -6 32 210
use FILL  FILL_37
timestamp 1018054153
transform 1 0 2864 0 -1 7680
box -16 -6 32 210
use FILL  FILL_38
timestamp 1018054153
transform 1 0 2880 0 -1 7680
box -16 -6 32 210
use FILL  FILL_39
timestamp 1018054153
transform 1 0 2896 0 -1 7680
box -16 -6 32 210
use FILL  FILL_40
timestamp 1018054153
transform 1 0 2912 0 -1 7680
box -16 -6 32 210
use FILL  FILL_41
timestamp 1018054153
transform 1 0 2928 0 -1 7680
box -16 -6 32 210
use FILL  FILL_42
timestamp 1018054153
transform 1 0 2944 0 -1 7680
box -16 -6 32 210
use FILL  FILL_43
timestamp 1018054153
transform 1 0 2960 0 -1 7680
box -16 -6 32 210
use FILL  FILL_44
timestamp 1018054153
transform 1 0 2976 0 -1 7680
box -16 -6 32 210
use FILL  FILL_45
timestamp 1018054153
transform 1 0 2992 0 -1 7680
box -16 -6 32 210
use FILL  FILL_46
timestamp 1018054153
transform 1 0 3008 0 -1 7680
box -16 -6 32 210
use FILL  FILL_47
timestamp 1018054153
transform 1 0 3024 0 -1 7680
box -16 -6 32 210
use FILL  FILL_48
timestamp 1018054153
transform 1 0 3040 0 -1 7680
box -16 -6 32 210
use FILL  FILL_49
timestamp 1018054153
transform 1 0 3056 0 -1 7680
box -16 -6 32 210
use FILL  FILL_50
timestamp 1018054153
transform 1 0 3072 0 -1 7680
box -16 -6 32 210
use FILL  FILL_51
timestamp 1018054153
transform 1 0 3088 0 -1 7680
box -16 -6 32 210
use FILL  FILL_52
timestamp 1018054153
transform 1 0 3104 0 -1 7680
box -16 -6 32 210
use FILL  FILL_53
timestamp 1018054153
transform 1 0 3120 0 -1 7680
box -16 -6 32 210
use FILL  FILL_54
timestamp 1018054153
transform 1 0 3136 0 -1 7680
box -16 -6 32 210
use FILL  FILL_55
timestamp 1018054153
transform 1 0 3152 0 -1 7680
box -16 -6 32 210
use FILL  FILL_56
timestamp 1018054153
transform 1 0 3168 0 -1 7680
box -16 -6 32 210
use FILL  FILL_57
timestamp 1018054153
transform 1 0 3184 0 -1 7680
box -16 -6 32 210
use FILL  FILL_58
timestamp 1018054153
transform 1 0 3200 0 -1 7680
box -16 -6 32 210
use FILL  FILL_59
timestamp 1018054153
transform 1 0 3216 0 -1 7680
box -16 -6 32 210
use FILL  FILL_60
timestamp 1018054153
transform 1 0 3232 0 -1 7680
box -16 -6 32 210
use FILL  FILL_61
timestamp 1018054153
transform 1 0 3248 0 -1 7680
box -16 -6 32 210
use FILL  FILL_62
timestamp 1018054153
transform 1 0 3264 0 -1 7680
box -16 -6 32 210
use FILL  FILL_63
timestamp 1018054153
transform 1 0 3280 0 -1 7680
box -16 -6 32 210
use FILL  FILL_64
timestamp 1018054153
transform 1 0 3296 0 -1 7680
box -16 -6 32 210
use FILL  FILL_65
timestamp 1018054153
transform 1 0 3312 0 -1 7680
box -16 -6 32 210
use FILL  FILL_66
timestamp 1018054153
transform 1 0 3328 0 -1 7680
box -16 -6 32 210
use FILL  FILL_67
timestamp 1018054153
transform 1 0 3344 0 -1 7680
box -16 -6 32 210
use FILL  FILL_68
timestamp 1018054153
transform 1 0 3360 0 -1 7680
box -16 -6 32 210
use FILL  FILL_69
timestamp 1018054153
transform 1 0 3376 0 -1 7680
box -16 -6 32 210
use FILL  FILL_70
timestamp 1018054153
transform 1 0 3392 0 -1 7680
box -16 -6 32 210
use FILL  FILL_71
timestamp 1018054153
transform 1 0 3408 0 -1 7680
box -16 -6 32 210
use FILL  FILL_72
timestamp 1018054153
transform 1 0 3424 0 -1 7680
box -16 -6 32 210
use FILL  FILL_73
timestamp 1018054153
transform 1 0 3440 0 -1 7680
box -16 -6 32 210
use FILL  FILL_74
timestamp 1018054153
transform 1 0 3456 0 -1 7680
box -16 -6 32 210
use FILL  FILL_75
timestamp 1018054153
transform 1 0 3472 0 -1 7680
box -16 -6 32 210
use FILL  FILL_76
timestamp 1018054153
transform 1 0 3488 0 -1 7680
box -16 -6 32 210
use FILL  FILL_77
timestamp 1018054153
transform 1 0 3504 0 -1 7680
box -16 -6 32 210
use FILL  FILL_78
timestamp 1018054153
transform 1 0 3520 0 -1 7680
box -16 -6 32 210
use FILL  FILL_79
timestamp 1018054153
transform 1 0 3536 0 -1 7680
box -16 -6 32 210
use FILL  FILL_80
timestamp 1018054153
transform 1 0 3552 0 -1 7680
box -16 -6 32 210
use FILL  FILL_81
timestamp 1018054153
transform 1 0 3568 0 -1 7680
box -16 -6 32 210
use FILL  FILL_82
timestamp 1018054153
transform 1 0 3584 0 -1 7680
box -16 -6 32 210
use FILL  FILL_83
timestamp 1018054153
transform 1 0 3600 0 -1 7680
box -16 -6 32 210
use FILL  FILL_84
timestamp 1018054153
transform 1 0 3616 0 -1 7680
box -16 -6 32 210
use FILL  FILL_85
timestamp 1018054153
transform 1 0 3632 0 -1 7680
box -16 -6 32 210
use FILL  FILL_86
timestamp 1018054153
transform 1 0 3648 0 -1 7680
box -16 -6 32 210
use FILL  FILL_87
timestamp 1018054153
transform 1 0 3664 0 -1 7680
box -16 -6 32 210
use FILL  FILL_88
timestamp 1018054153
transform 1 0 3680 0 -1 7680
box -16 -6 32 210
use FILL  FILL_89
timestamp 1018054153
transform 1 0 3696 0 -1 7680
box -16 -6 32 210
use FILL  FILL_90
timestamp 1018054153
transform 1 0 3712 0 -1 7680
box -16 -6 32 210
use FILL  FILL_91
timestamp 1018054153
transform 1 0 3728 0 -1 7680
box -16 -6 32 210
use FILL  FILL_92
timestamp 1018054153
transform 1 0 3744 0 -1 7680
box -16 -6 32 210
use FILL  FILL_93
timestamp 1018054153
transform 1 0 3760 0 -1 7680
box -16 -6 32 210
use FILL  FILL_94
timestamp 1018054153
transform 1 0 3776 0 -1 7680
box -16 -6 32 210
use FILL  FILL_95
timestamp 1018054153
transform 1 0 3792 0 -1 7680
box -16 -6 32 210
use FILL  FILL_96
timestamp 1018054153
transform 1 0 3808 0 -1 7680
box -16 -6 32 210
use FILL  FILL_97
timestamp 1018054153
transform 1 0 3824 0 -1 7680
box -16 -6 32 210
use FILL  FILL_98
timestamp 1018054153
transform 1 0 3840 0 -1 7680
box -16 -6 32 210
use FILL  FILL_99
timestamp 1018054153
transform 1 0 3856 0 -1 7680
box -16 -6 32 210
use FILL  FILL_100
timestamp 1018054153
transform 1 0 3872 0 -1 7680
box -16 -6 32 210
use FILL  FILL_101
timestamp 1018054153
transform 1 0 3888 0 -1 7680
box -16 -6 32 210
use FILL  FILL_102
timestamp 1018054153
transform 1 0 3904 0 -1 7680
box -16 -6 32 210
use FILL  FILL_103
timestamp 1018054153
transform 1 0 3920 0 -1 7680
box -16 -6 32 210
use FILL  FILL_104
timestamp 1018054153
transform 1 0 3936 0 -1 7680
box -16 -6 32 210
use FILL  FILL_105
timestamp 1018054153
transform 1 0 3952 0 -1 7680
box -16 -6 32 210
use FILL  FILL_106
timestamp 1018054153
transform 1 0 3968 0 -1 7680
box -16 -6 32 210
use FILL  FILL_107
timestamp 1018054153
transform 1 0 3984 0 -1 7680
box -16 -6 32 210
use FILL  FILL_108
timestamp 1018054153
transform 1 0 4000 0 -1 7680
box -16 -6 32 210
use FILL  FILL_109
timestamp 1018054153
transform 1 0 4016 0 -1 7680
box -16 -6 32 210
use FILL  FILL_110
timestamp 1018054153
transform 1 0 4032 0 -1 7680
box -16 -6 32 210
use FILL  FILL_111
timestamp 1018054153
transform 1 0 4048 0 -1 7680
box -16 -6 32 210
use FILL  FILL_112
timestamp 1018054153
transform 1 0 4064 0 -1 7680
box -16 -6 32 210
use FILL  FILL_113
timestamp 1018054153
transform 1 0 4080 0 -1 7680
box -16 -6 32 210
use FILL  FILL_114
timestamp 1018054153
transform 1 0 4096 0 -1 7680
box -16 -6 32 210
use FILL  FILL_115
timestamp 1018054153
transform 1 0 4112 0 -1 7680
box -16 -6 32 210
use FILL  FILL_116
timestamp 1018054153
transform 1 0 4128 0 -1 7680
box -16 -6 32 210
use FILL  FILL_117
timestamp 1018054153
transform 1 0 4144 0 -1 7680
box -16 -6 32 210
use FILL  FILL_118
timestamp 1018054153
transform 1 0 4160 0 -1 7680
box -16 -6 32 210
use FILL  FILL_119
timestamp 1018054153
transform 1 0 4176 0 -1 7680
box -16 -6 32 210
use FILL  FILL_120
timestamp 1018054153
transform 1 0 4192 0 -1 7680
box -16 -6 32 210
use FILL  FILL_121
timestamp 1018054153
transform 1 0 4208 0 -1 7680
box -16 -6 32 210
use FILL  FILL_122
timestamp 1018054153
transform 1 0 4224 0 -1 7680
box -16 -6 32 210
use FILL  FILL_123
timestamp 1018054153
transform 1 0 4240 0 -1 7680
box -16 -6 32 210
use FILL  FILL_124
timestamp 1018054153
transform 1 0 4256 0 -1 7680
box -16 -6 32 210
use FILL  FILL_125
timestamp 1018054153
transform 1 0 4272 0 -1 7680
box -16 -6 32 210
use FILL  FILL_126
timestamp 1018054153
transform 1 0 4288 0 -1 7680
box -16 -6 32 210
use FILL  FILL_127
timestamp 1018054153
transform 1 0 4304 0 -1 7680
box -16 -6 32 210
use FILL  FILL_128
timestamp 1018054153
transform 1 0 4320 0 -1 7680
box -16 -6 32 210
use FILL  FILL_129
timestamp 1018054153
transform 1 0 4336 0 -1 7680
box -16 -6 32 210
use FILL  FILL_130
timestamp 1018054153
transform 1 0 4352 0 -1 7680
box -16 -6 32 210
use FILL  FILL_131
timestamp 1018054153
transform 1 0 4368 0 -1 7680
box -16 -6 32 210
use FILL  FILL_132
timestamp 1018054153
transform 1 0 4384 0 -1 7680
box -16 -6 32 210
use FILL  FILL_133
timestamp 1018054153
transform 1 0 4400 0 -1 7680
box -16 -6 32 210
use FILL  FILL_134
timestamp 1018054153
transform 1 0 4416 0 -1 7680
box -16 -6 32 210
use FILL  FILL_135
timestamp 1018054153
transform 1 0 4432 0 -1 7680
box -16 -6 32 210
use FILL  FILL_136
timestamp 1018054153
transform 1 0 4448 0 -1 7680
box -16 -6 32 210
use FILL  FILL_137
timestamp 1018054153
transform 1 0 4464 0 -1 7680
box -16 -6 32 210
use FILL  FILL_138
timestamp 1018054153
transform 1 0 4480 0 -1 7680
box -16 -6 32 210
use FILL  FILL_139
timestamp 1018054153
transform 1 0 4496 0 -1 7680
box -16 -6 32 210
use FILL  FILL_140
timestamp 1018054153
transform 1 0 4512 0 -1 7680
box -16 -6 32 210
use FILL  FILL_141
timestamp 1018054153
transform 1 0 4528 0 -1 7680
box -16 -6 32 210
use FILL  FILL_142
timestamp 1018054153
transform 1 0 4544 0 -1 7680
box -16 -6 32 210
use FILL  FILL_143
timestamp 1018054153
transform 1 0 4560 0 -1 7680
box -16 -6 32 210
use FILL  FILL_144
timestamp 1018054153
transform 1 0 4576 0 -1 7680
box -16 -6 32 210
use FILL  FILL_145
timestamp 1018054153
transform 1 0 4592 0 -1 7680
box -16 -6 32 210
use FILL  FILL_146
timestamp 1018054153
transform 1 0 4608 0 -1 7680
box -16 -6 32 210
use FILL  FILL_147
timestamp 1018054153
transform 1 0 4624 0 -1 7680
box -16 -6 32 210
use FILL  FILL_148
timestamp 1018054153
transform 1 0 4640 0 -1 7680
box -16 -6 32 210
use FILL  FILL_149
timestamp 1018054153
transform 1 0 4656 0 -1 7680
box -16 -6 32 210
use FILL  FILL_150
timestamp 1018054153
transform 1 0 4672 0 -1 7680
box -16 -6 32 210
use FILL  FILL_151
timestamp 1018054153
transform 1 0 4688 0 -1 7680
box -16 -6 32 210
use FILL  FILL_152
timestamp 1018054153
transform 1 0 4704 0 -1 7680
box -16 -6 32 210
use FILL  FILL_153
timestamp 1018054153
transform 1 0 4720 0 -1 7680
box -16 -6 32 210
use FILL  FILL_154
timestamp 1018054153
transform 1 0 4736 0 -1 7680
box -16 -6 32 210
use FILL  FILL_155
timestamp 1018054153
transform 1 0 4752 0 -1 7680
box -16 -6 32 210
use FILL  FILL_156
timestamp 1018054153
transform 1 0 4768 0 -1 7680
box -16 -6 32 210
use FILL  FILL_157
timestamp 1018054153
transform 1 0 4784 0 -1 7680
box -16 -6 32 210
use FILL  FILL_158
timestamp 1018054153
transform 1 0 4800 0 -1 7680
box -16 -6 32 210
use FILL  FILL_159
timestamp 1018054153
transform 1 0 4816 0 -1 7680
box -16 -6 32 210
use FILL  FILL_160
timestamp 1018054153
transform 1 0 4832 0 -1 7680
box -16 -6 32 210
use FILL  FILL_161
timestamp 1018054153
transform 1 0 4848 0 -1 7680
box -16 -6 32 210
use FILL  FILL_162
timestamp 1018054153
transform 1 0 4864 0 -1 7680
box -16 -6 32 210
use FILL  FILL_163
timestamp 1018054153
transform 1 0 4880 0 -1 7680
box -16 -6 32 210
use FILL  FILL_164
timestamp 1018054153
transform 1 0 4896 0 -1 7680
box -16 -6 32 210
use FILL  FILL_165
timestamp 1018054153
transform 1 0 4912 0 -1 7680
box -16 -6 32 210
use FILL  FILL_166
timestamp 1018054153
transform 1 0 4928 0 -1 7680
box -16 -6 32 210
use FILL  FILL_167
timestamp 1018054153
transform 1 0 4944 0 -1 7680
box -16 -6 32 210
use FILL  FILL_168
timestamp 1018054153
transform 1 0 4960 0 -1 7680
box -16 -6 32 210
use FILL  FILL_169
timestamp 1018054153
transform 1 0 4976 0 -1 7680
box -16 -6 32 210
use FILL  FILL_170
timestamp 1018054153
transform 1 0 4992 0 -1 7680
box -16 -6 32 210
use FILL  FILL_171
timestamp 1018054153
transform 1 0 5008 0 -1 7680
box -16 -6 32 210
use FILL  FILL_172
timestamp 1018054153
transform 1 0 5024 0 -1 7680
box -16 -6 32 210
use FILL  FILL_173
timestamp 1018054153
transform 1 0 5040 0 -1 7680
box -16 -6 32 210
use FILL  FILL_174
timestamp 1018054153
transform 1 0 5056 0 -1 7680
box -16 -6 32 210
use FILL  FILL_175
timestamp 1018054153
transform 1 0 5072 0 -1 7680
box -16 -6 32 210
use FILL  FILL_176
timestamp 1018054153
transform 1 0 5088 0 -1 7680
box -16 -6 32 210
use FILL  FILL_177
timestamp 1018054153
transform 1 0 5104 0 -1 7680
box -16 -6 32 210
use FILL  FILL_178
timestamp 1018054153
transform 1 0 5120 0 -1 7680
box -16 -6 32 210
use FILL  FILL_179
timestamp 1018054153
transform 1 0 5136 0 -1 7680
box -16 -6 32 210
use FILL  FILL_180
timestamp 1018054153
transform 1 0 5152 0 -1 7680
box -16 -6 32 210
use FILL  FILL_181
timestamp 1018054153
transform 1 0 5168 0 -1 7680
box -16 -6 32 210
use FILL  FILL_182
timestamp 1018054153
transform 1 0 5184 0 -1 7680
box -16 -6 32 210
use FILL  FILL_183
timestamp 1018054153
transform 1 0 5200 0 -1 7680
box -16 -6 32 210
use FILL  FILL_184
timestamp 1018054153
transform 1 0 5216 0 -1 7680
box -16 -6 32 210
use FILL  FILL_185
timestamp 1018054153
transform 1 0 5232 0 -1 7680
box -16 -6 32 210
use FILL  FILL_186
timestamp 1018054153
transform 1 0 5248 0 -1 7680
box -16 -6 32 210
use FILL  FILL_187
timestamp 1018054153
transform 1 0 5264 0 -1 7680
box -16 -6 32 210
use FILL  FILL_188
timestamp 1018054153
transform 1 0 5280 0 -1 7680
box -16 -6 32 210
use FILL  FILL_189
timestamp 1018054153
transform 1 0 5296 0 -1 7680
box -16 -6 32 210
use FILL  FILL_190
timestamp 1018054153
transform 1 0 5312 0 -1 7680
box -16 -6 32 210
use FILL  FILL_191
timestamp 1018054153
transform 1 0 5328 0 -1 7680
box -16 -6 32 210
use FILL  FILL_192
timestamp 1018054153
transform 1 0 5344 0 -1 7680
box -16 -6 32 210
use FILL  FILL_193
timestamp 1018054153
transform 1 0 5360 0 -1 7680
box -16 -6 32 210
use FILL  FILL_194
timestamp 1018054153
transform 1 0 5376 0 -1 7680
box -16 -6 32 210
use FILL  FILL_195
timestamp 1018054153
transform 1 0 5392 0 -1 7680
box -16 -6 32 210
use FILL  FILL_196
timestamp 1018054153
transform 1 0 5408 0 -1 7680
box -16 -6 32 210
use FILL  FILL_197
timestamp 1018054153
transform 1 0 5424 0 -1 7680
box -16 -6 32 210
use FILL  FILL_198
timestamp 1018054153
transform 1 0 5440 0 -1 7680
box -16 -6 32 210
use FILL  FILL_199
timestamp 1018054153
transform 1 0 5456 0 -1 7680
box -16 -6 32 210
use FILL  FILL_200
timestamp 1018054153
transform 1 0 5472 0 -1 7680
box -16 -6 32 210
use FILL  FILL_201
timestamp 1018054153
transform 1 0 5488 0 -1 7680
box -16 -6 32 210
use FILL  FILL_202
timestamp 1018054153
transform 1 0 5504 0 -1 7680
box -16 -6 32 210
use FILL  FILL_203
timestamp 1018054153
transform 1 0 5520 0 -1 7680
box -16 -6 32 210
use FILL  FILL_204
timestamp 1018054153
transform 1 0 5536 0 -1 7680
box -16 -6 32 210
use FILL  FILL_205
timestamp 1018054153
transform 1 0 5552 0 -1 7680
box -16 -6 32 210
use FILL  FILL_206
timestamp 1018054153
transform 1 0 5568 0 -1 7680
box -16 -6 32 210
use FILL  FILL_207
timestamp 1018054153
transform 1 0 5584 0 -1 7680
box -16 -6 32 210
use FILL  FILL_208
timestamp 1018054153
transform 1 0 5600 0 -1 7680
box -16 -6 32 210
use FILL  FILL_209
timestamp 1018054153
transform 1 0 5616 0 -1 7680
box -16 -6 32 210
use FILL  FILL_210
timestamp 1018054153
transform 1 0 5632 0 -1 7680
box -16 -6 32 210
use FILL  FILL_211
timestamp 1018054153
transform 1 0 5648 0 -1 7680
box -16 -6 32 210
use FILL  FILL_212
timestamp 1018054153
transform 1 0 5664 0 -1 7680
box -16 -6 32 210
use FILL  FILL_213
timestamp 1018054153
transform 1 0 5680 0 -1 7680
box -16 -6 32 210
use FILL  FILL_214
timestamp 1018054153
transform 1 0 5696 0 -1 7680
box -16 -6 32 210
use FILL  FILL_215
timestamp 1018054153
transform 1 0 5712 0 -1 7680
box -16 -6 32 210
use FILL  FILL_216
timestamp 1018054153
transform 1 0 5728 0 -1 7680
box -16 -6 32 210
use FILL  FILL_217
timestamp 1018054153
transform 1 0 5744 0 -1 7680
box -16 -6 32 210
use FILL  FILL_218
timestamp 1018054153
transform 1 0 5760 0 -1 7680
box -16 -6 32 210
use FILL  FILL_219
timestamp 1018054153
transform 1 0 5776 0 -1 7680
box -16 -6 32 210
use FILL  FILL_220
timestamp 1018054153
transform 1 0 5792 0 -1 7680
box -16 -6 32 210
use FILL  FILL_221
timestamp 1018054153
transform 1 0 5808 0 -1 7680
box -16 -6 32 210
use FILL  FILL_222
timestamp 1018054153
transform 1 0 5824 0 -1 7680
box -16 -6 32 210
use FILL  FILL_223
timestamp 1018054153
transform 1 0 5840 0 -1 7680
box -16 -6 32 210
use FILL  FILL_224
timestamp 1018054153
transform 1 0 5856 0 -1 7680
box -16 -6 32 210
use FILL  FILL_225
timestamp 1018054153
transform 1 0 5872 0 -1 7680
box -16 -6 32 210
use FILL  FILL_226
timestamp 1018054153
transform 1 0 5888 0 -1 7680
box -16 -6 32 210
use FILL  FILL_227
timestamp 1018054153
transform 1 0 5904 0 -1 7680
box -16 -6 32 210
use FILL  FILL_228
timestamp 1018054153
transform 1 0 5920 0 -1 7680
box -16 -6 32 210
use FILL  FILL_229
timestamp 1018054153
transform 1 0 5936 0 -1 7680
box -16 -6 32 210
use FILL  FILL_230
timestamp 1018054153
transform 1 0 5952 0 -1 7680
box -16 -6 32 210
use FILL  FILL_231
timestamp 1018054153
transform 1 0 5968 0 -1 7680
box -16 -6 32 210
use FILL  FILL_232
timestamp 1018054153
transform 1 0 5984 0 -1 7680
box -16 -6 32 210
use FILL  FILL_233
timestamp 1018054153
transform 1 0 6000 0 -1 7680
box -16 -6 32 210
use FILL  FILL_234
timestamp 1018054153
transform 1 0 6016 0 -1 7680
box -16 -6 32 210
use FILL  FILL_235
timestamp 1018054153
transform 1 0 6032 0 -1 7680
box -16 -6 32 210
use FILL  FILL_236
timestamp 1018054153
transform 1 0 6048 0 -1 7680
box -16 -6 32 210
use FILL  FILL_237
timestamp 1018054153
transform 1 0 6064 0 -1 7680
box -16 -6 32 210
use FILL  FILL_238
timestamp 1018054153
transform 1 0 6080 0 -1 7680
box -16 -6 32 210
use FILL  FILL_239
timestamp 1018054153
transform 1 0 6096 0 -1 7680
box -16 -6 32 210
use FILL  FILL_240
timestamp 1018054153
transform 1 0 6112 0 -1 7680
box -16 -6 32 210
use FILL  FILL_241
timestamp 1018054153
transform 1 0 6128 0 -1 7680
box -16 -6 32 210
use FILL  FILL_242
timestamp 1018054153
transform 1 0 6144 0 -1 7680
box -16 -6 32 210
use FILL  FILL_243
timestamp 1018054153
transform 1 0 6160 0 -1 7680
box -16 -6 32 210
use FILL  FILL_244
timestamp 1018054153
transform 1 0 6176 0 -1 7680
box -16 -6 32 210
use FILL  FILL_245
timestamp 1018054153
transform 1 0 6192 0 -1 7680
box -16 -6 32 210
use FILL  FILL_246
timestamp 1018054153
transform 1 0 6208 0 -1 7680
box -16 -6 32 210
use FILL  FILL_247
timestamp 1018054153
transform 1 0 6224 0 -1 7680
box -16 -6 32 210
use FILL  FILL_248
timestamp 1018054153
transform 1 0 6240 0 -1 7680
box -16 -6 32 210
use FILL  FILL_249
timestamp 1018054153
transform 1 0 6256 0 -1 7680
box -16 -6 32 210
use FILL  FILL_250
timestamp 1018054153
transform 1 0 6272 0 -1 7680
box -16 -6 32 210
use FILL  FILL_251
timestamp 1018054153
transform 1 0 6288 0 -1 7680
box -16 -6 32 210
use FILL  FILL_252
timestamp 1018054153
transform 1 0 6304 0 -1 7680
box -16 -6 32 210
use FILL  FILL_253
timestamp 1018054153
transform 1 0 6320 0 -1 7680
box -16 -6 32 210
use FILL  FILL_254
timestamp 1018054153
transform 1 0 6336 0 -1 7680
box -16 -6 32 210
use FILL  FILL_255
timestamp 1018054153
transform 1 0 6352 0 -1 7680
box -16 -6 32 210
use FILL  FILL_256
timestamp 1018054153
transform 1 0 6368 0 -1 7680
box -16 -6 32 210
use FILL  FILL_257
timestamp 1018054153
transform 1 0 6384 0 -1 7680
box -16 -6 32 210
use FILL  FILL_258
timestamp 1018054153
transform 1 0 6400 0 -1 7680
box -16 -6 32 210
use FILL  FILL_259
timestamp 1018054153
transform 1 0 6416 0 -1 7680
box -16 -6 32 210
use FILL  FILL_260
timestamp 1018054153
transform 1 0 6432 0 -1 7680
box -16 -6 32 210
use FILL  FILL_261
timestamp 1018054153
transform 1 0 6448 0 -1 7680
box -16 -6 32 210
use FILL  FILL_262
timestamp 1018054153
transform 1 0 6464 0 -1 7680
box -16 -6 32 210
use FILL  FILL_263
timestamp 1018054153
transform 1 0 6480 0 -1 7680
box -16 -6 32 210
use FILL  FILL_264
timestamp 1018054153
transform 1 0 6496 0 -1 7680
box -16 -6 32 210
use FILL  FILL_265
timestamp 1018054153
transform 1 0 6512 0 -1 7680
box -16 -6 32 210
use FILL  FILL_266
timestamp 1018054153
transform 1 0 6528 0 -1 7680
box -16 -6 32 210
use FILL  FILL_267
timestamp 1018054153
transform 1 0 6544 0 -1 7680
box -16 -6 32 210
use FILL  FILL_268
timestamp 1018054153
transform 1 0 6560 0 -1 7680
box -16 -6 32 210
use FILL  FILL_269
timestamp 1018054153
transform 1 0 6576 0 -1 7680
box -16 -6 32 210
use FILL  FILL_270
timestamp 1018054153
transform 1 0 6592 0 -1 7680
box -16 -6 32 210
use FILL  FILL_271
timestamp 1018054153
transform 1 0 6608 0 -1 7680
box -16 -6 32 210
use FILL  FILL_272
timestamp 1018054153
transform 1 0 6624 0 -1 7680
box -16 -6 32 210
use FILL  FILL_273
timestamp 1018054153
transform 1 0 6640 0 -1 7680
box -16 -6 32 210
use FILL  FILL_274
timestamp 1018054153
transform 1 0 6656 0 -1 7680
box -16 -6 32 210
use FILL  FILL_275
timestamp 1018054153
transform 1 0 6672 0 -1 7680
box -16 -6 32 210
use FILL  FILL_276
timestamp 1018054153
transform 1 0 6688 0 -1 7680
box -16 -6 32 210
use FILL  FILL_277
timestamp 1018054153
transform 1 0 6704 0 -1 7680
box -16 -6 32 210
use FILL  FILL_278
timestamp 1018054153
transform 1 0 6720 0 -1 7680
box -16 -6 32 210
use FILL  FILL_279
timestamp 1018054153
transform 1 0 6736 0 -1 7680
box -16 -6 32 210
use FILL  FILL_280
timestamp 1018054153
transform 1 0 6752 0 -1 7680
box -16 -6 32 210
use FILL  FILL_281
timestamp 1018054153
transform 1 0 6768 0 -1 7680
box -16 -6 32 210
use FILL  FILL_282
timestamp 1018054153
transform 1 0 6784 0 -1 7680
box -16 -6 32 210
use FILL  FILL_283
timestamp 1018054153
transform 1 0 6800 0 -1 7680
box -16 -6 32 210
use FILL  FILL_284
timestamp 1018054153
transform 1 0 6816 0 -1 7680
box -16 -6 32 210
use FILL  FILL_285
timestamp 1018054153
transform 1 0 6832 0 -1 7680
box -16 -6 32 210
use FILL  FILL_286
timestamp 1018054153
transform 1 0 6848 0 -1 7680
box -16 -6 32 210
use FILL  FILL_287
timestamp 1018054153
transform 1 0 6864 0 -1 7680
box -16 -6 32 210
use FILL  FILL_288
timestamp 1018054153
transform 1 0 6880 0 -1 7680
box -16 -6 32 210
use FILL  FILL_289
timestamp 1018054153
transform 1 0 6896 0 -1 7680
box -16 -6 32 210
use FILL  FILL_290
timestamp 1018054153
transform 1 0 6912 0 -1 7680
box -16 -6 32 210
use FILL  FILL_291
timestamp 1018054153
transform 1 0 6928 0 -1 7680
box -16 -6 32 210
use FILL  FILL_292
timestamp 1018054153
transform 1 0 6944 0 -1 7680
box -16 -6 32 210
use FILL  FILL_293
timestamp 1018054153
transform 1 0 6960 0 -1 7680
box -16 -6 32 210
use FILL  FILL_294
timestamp 1018054153
transform 1 0 6976 0 -1 7680
box -16 -6 32 210
use FILL  FILL_295
timestamp 1018054153
transform 1 0 6992 0 -1 7680
box -16 -6 32 210
use FILL  FILL_296
timestamp 1018054153
transform 1 0 7008 0 -1 7680
box -16 -6 32 210
use FILL  FILL_297
timestamp 1018054153
transform 1 0 7024 0 -1 7680
box -16 -6 32 210
use FILL  FILL_298
timestamp 1018054153
transform 1 0 7040 0 -1 7680
box -16 -6 32 210
use FILL  FILL_299
timestamp 1018054153
transform 1 0 7056 0 -1 7680
box -16 -6 32 210
use FILL  FILL_300
timestamp 1018054153
transform 1 0 7072 0 -1 7680
box -16 -6 32 210
use FILL  FILL_301
timestamp 1018054153
transform 1 0 7088 0 -1 7680
box -16 -6 32 210
use FILL  FILL_302
timestamp 1018054153
transform 1 0 7104 0 -1 7680
box -16 -6 32 210
use FILL  FILL_303
timestamp 1018054153
transform 1 0 7120 0 -1 7680
box -16 -6 32 210
use FILL  FILL_304
timestamp 1018054153
transform 1 0 7136 0 -1 7680
box -16 -6 32 210
use FILL  FILL_305
timestamp 1018054153
transform 1 0 7152 0 -1 7680
box -16 -6 32 210
use FILL  FILL_306
timestamp 1018054153
transform 1 0 7168 0 -1 7680
box -16 -6 32 210
use FILL  FILL_307
timestamp 1018054153
transform 1 0 7184 0 -1 7680
box -16 -6 32 210
use FILL  FILL_308
timestamp 1018054153
transform 1 0 7200 0 -1 7680
box -16 -6 32 210
use FILL  FILL_309
timestamp 1018054153
transform 1 0 7216 0 -1 7680
box -16 -6 32 210
use FILL  FILL_310
timestamp 1018054153
transform 1 0 7232 0 -1 7680
box -16 -6 32 210
use FILL  FILL_311
timestamp 1018054153
transform 1 0 7248 0 -1 7680
box -16 -6 32 210
use FILL  FILL_312
timestamp 1018054153
transform 1 0 7264 0 -1 7680
box -16 -6 32 210
use FILL  FILL_313
timestamp 1018054153
transform 1 0 7280 0 -1 7680
box -16 -6 32 210
use FILL  FILL_314
timestamp 1018054153
transform 1 0 7296 0 -1 7680
box -16 -6 32 210
use FILL  FILL_315
timestamp 1018054153
transform 1 0 7312 0 -1 7680
box -16 -6 32 210
use FILL  FILL_316
timestamp 1018054153
transform 1 0 7328 0 -1 7680
box -16 -6 32 210
use FILL  FILL_317
timestamp 1018054153
transform 1 0 7344 0 -1 7680
box -16 -6 32 210
use FILL  FILL_318
timestamp 1018054153
transform 1 0 7360 0 -1 7680
box -16 -6 32 210
use FILL  FILL_319
timestamp 1018054153
transform 1 0 7376 0 -1 7680
box -16 -6 32 210
use FILL  FILL_320
timestamp 1018054153
transform 1 0 7392 0 -1 7680
box -16 -6 32 210
use FILL  FILL_321
timestamp 1018054153
transform 1 0 7408 0 -1 7680
box -16 -6 32 210
use FILL  FILL_322
timestamp 1018054153
transform 1 0 7424 0 -1 7680
box -16 -6 32 210
use FILL  FILL_323
timestamp 1018054153
transform 1 0 7440 0 -1 7680
box -16 -6 32 210
use FILL  FILL_324
timestamp 1018054153
transform 1 0 7456 0 -1 7680
box -16 -6 32 210
use FILL  FILL_325
timestamp 1018054153
transform 1 0 7472 0 -1 7680
box -16 -6 32 210
use FILL  FILL_326
timestamp 1018054153
transform 1 0 7488 0 -1 7680
box -16 -6 32 210
use FILL  FILL_327
timestamp 1018054153
transform 1 0 7504 0 -1 7680
box -16 -6 32 210
use FILL  FILL_328
timestamp 1018054153
transform 1 0 7520 0 -1 7680
box -16 -6 32 210
use FILL  FILL_329
timestamp 1018054153
transform 1 0 7536 0 -1 7680
box -16 -6 32 210
use FILL  FILL_330
timestamp 1018054153
transform 1 0 7552 0 -1 7680
box -16 -6 32 210
use FILL  FILL_331
timestamp 1018054153
transform 1 0 7568 0 -1 7680
box -16 -6 32 210
use FILL  FILL_332
timestamp 1018054153
transform 1 0 7584 0 -1 7680
box -16 -6 32 210
use FILL  FILL_333
timestamp 1018054153
transform 1 0 7600 0 -1 7680
box -16 -6 32 210
use FILL  FILL_334
timestamp 1018054153
transform 1 0 7616 0 -1 7680
box -16 -6 32 210
use FILL  FILL_335
timestamp 1018054153
transform 1 0 7632 0 -1 7680
box -16 -6 32 210
use FILL  FILL_336
timestamp 1018054153
transform 1 0 7648 0 -1 7680
box -16 -6 32 210
use FILL  FILL_337
timestamp 1018054153
transform 1 0 7664 0 -1 7680
box -16 -6 32 210
use FILL  FILL_338
timestamp 1018054153
transform 1 0 7680 0 -1 7680
box -16 -6 32 210
use FILL  FILL_339
timestamp 1018054153
transform 1 0 7696 0 -1 7680
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_1
timestamp 1542725905
transform 1 0 7788 0 1 7480
box -48 -6 48 6
use FILL  FILL_340
timestamp 1018054153
transform 1 0 7712 0 -1 7680
box -16 -6 32 210
use M2_M1  M2_M1_0
timestamp 1542725905
transform 1 0 4456 0 1 7410
box -4 -4 4 4
use M2_M1  M2_M1_1
timestamp 1542725905
transform 1 0 5528 0 1 7410
box -4 -4 4 4
use PADGND  PADGND_0
timestamp 1084294269
transform 0 1 8000 -1 0 8000
box -6 -6 606 2000
use mult_pad_VIA1  mult_pad_VIA1_2
timestamp 1542725905
transform 1 0 2092 0 1 7280
box -48 -6 48 6
use FILL  FILL_341
timestamp 1018054153
transform 1 0 2272 0 1 7280
box -16 -6 32 210
use FILL  FILL_343
timestamp 1018054153
transform 1 0 2288 0 1 7280
box -16 -6 32 210
use FILL  FILL_345
timestamp 1018054153
transform 1 0 2304 0 1 7280
box -16 -6 32 210
use FILL  FILL_347
timestamp 1018054153
transform 1 0 2320 0 1 7280
box -16 -6 32 210
use FILL  FILL_349
timestamp 1018054153
transform 1 0 2336 0 1 7280
box -16 -6 32 210
use FILL  FILL_351
timestamp 1018054153
transform 1 0 2352 0 1 7280
box -16 -6 32 210
use FILL  FILL_353
timestamp 1018054153
transform 1 0 2368 0 1 7280
box -16 -6 32 210
use FILL  FILL_355
timestamp 1018054153
transform 1 0 2384 0 1 7280
box -16 -6 32 210
use FILL  FILL_357
timestamp 1018054153
transform 1 0 2400 0 1 7280
box -16 -6 32 210
use FILL  FILL_359
timestamp 1018054153
transform 1 0 2416 0 1 7280
box -16 -6 32 210
use FILL  FILL_361
timestamp 1018054153
transform 1 0 2432 0 1 7280
box -16 -6 32 210
use FILL  FILL_363
timestamp 1018054153
transform 1 0 2448 0 1 7280
box -16 -6 32 210
use FILL  FILL_365
timestamp 1018054153
transform 1 0 2464 0 1 7280
box -16 -6 32 210
use FILL  FILL_367
timestamp 1018054153
transform 1 0 2480 0 1 7280
box -16 -6 32 210
use FILL  FILL_369
timestamp 1018054153
transform 1 0 2496 0 1 7280
box -16 -6 32 210
use FILL  FILL_371
timestamp 1018054153
transform 1 0 2512 0 1 7280
box -16 -6 32 210
use FILL  FILL_373
timestamp 1018054153
transform 1 0 2528 0 1 7280
box -16 -6 32 210
use FILL  FILL_375
timestamp 1018054153
transform 1 0 2544 0 1 7280
box -16 -6 32 210
use FILL  FILL_377
timestamp 1018054153
transform 1 0 2560 0 1 7280
box -16 -6 32 210
use FILL  FILL_379
timestamp 1018054153
transform 1 0 2576 0 1 7280
box -16 -6 32 210
use FILL  FILL_381
timestamp 1018054153
transform 1 0 2592 0 1 7280
box -16 -6 32 210
use FILL  FILL_383
timestamp 1018054153
transform 1 0 2608 0 1 7280
box -16 -6 32 210
use FILL  FILL_385
timestamp 1018054153
transform 1 0 2624 0 1 7280
box -16 -6 32 210
use FILL  FILL_387
timestamp 1018054153
transform 1 0 2640 0 1 7280
box -16 -6 32 210
use FILL  FILL_389
timestamp 1018054153
transform 1 0 2656 0 1 7280
box -16 -6 32 210
use FILL  FILL_391
timestamp 1018054153
transform 1 0 2672 0 1 7280
box -16 -6 32 210
use FILL  FILL_393
timestamp 1018054153
transform 1 0 2688 0 1 7280
box -16 -6 32 210
use FILL  FILL_395
timestamp 1018054153
transform 1 0 2704 0 1 7280
box -16 -6 32 210
use FILL  FILL_397
timestamp 1018054153
transform 1 0 2720 0 1 7280
box -16 -6 32 210
use FILL  FILL_399
timestamp 1018054153
transform 1 0 2736 0 1 7280
box -16 -6 32 210
use FILL  FILL_401
timestamp 1018054153
transform 1 0 2752 0 1 7280
box -16 -6 32 210
use FILL  FILL_403
timestamp 1018054153
transform 1 0 2768 0 1 7280
box -16 -6 32 210
use FILL  FILL_405
timestamp 1018054153
transform 1 0 2784 0 1 7280
box -16 -6 32 210
use FILL  FILL_407
timestamp 1018054153
transform 1 0 2800 0 1 7280
box -16 -6 32 210
use FILL  FILL_409
timestamp 1018054153
transform 1 0 2816 0 1 7280
box -16 -6 32 210
use FILL  FILL_411
timestamp 1018054153
transform 1 0 2832 0 1 7280
box -16 -6 32 210
use FILL  FILL_413
timestamp 1018054153
transform 1 0 2848 0 1 7280
box -16 -6 32 210
use FILL  FILL_415
timestamp 1018054153
transform 1 0 2864 0 1 7280
box -16 -6 32 210
use FILL  FILL_417
timestamp 1018054153
transform 1 0 2880 0 1 7280
box -16 -6 32 210
use FILL  FILL_419
timestamp 1018054153
transform 1 0 2896 0 1 7280
box -16 -6 32 210
use FILL  FILL_421
timestamp 1018054153
transform 1 0 2912 0 1 7280
box -16 -6 32 210
use FILL  FILL_423
timestamp 1018054153
transform 1 0 2928 0 1 7280
box -16 -6 32 210
use FILL  FILL_425
timestamp 1018054153
transform 1 0 2944 0 1 7280
box -16 -6 32 210
use FILL  FILL_427
timestamp 1018054153
transform 1 0 2960 0 1 7280
box -16 -6 32 210
use FILL  FILL_429
timestamp 1018054153
transform 1 0 2976 0 1 7280
box -16 -6 32 210
use FILL  FILL_431
timestamp 1018054153
transform 1 0 2992 0 1 7280
box -16 -6 32 210
use FILL  FILL_433
timestamp 1018054153
transform 1 0 3008 0 1 7280
box -16 -6 32 210
use FILL  FILL_435
timestamp 1018054153
transform 1 0 3024 0 1 7280
box -16 -6 32 210
use FILL  FILL_437
timestamp 1018054153
transform 1 0 3040 0 1 7280
box -16 -6 32 210
use FILL  FILL_439
timestamp 1018054153
transform 1 0 3056 0 1 7280
box -16 -6 32 210
use FILL  FILL_441
timestamp 1018054153
transform 1 0 3072 0 1 7280
box -16 -6 32 210
use FILL  FILL_443
timestamp 1018054153
transform 1 0 3088 0 1 7280
box -16 -6 32 210
use FILL  FILL_445
timestamp 1018054153
transform 1 0 3104 0 1 7280
box -16 -6 32 210
use FILL  FILL_447
timestamp 1018054153
transform 1 0 3120 0 1 7280
box -16 -6 32 210
use FILL  FILL_449
timestamp 1018054153
transform 1 0 3136 0 1 7280
box -16 -6 32 210
use FILL  FILL_451
timestamp 1018054153
transform 1 0 3152 0 1 7280
box -16 -6 32 210
use FILL  FILL_453
timestamp 1018054153
transform 1 0 3168 0 1 7280
box -16 -6 32 210
use FILL  FILL_455
timestamp 1018054153
transform 1 0 3184 0 1 7280
box -16 -6 32 210
use FILL  FILL_457
timestamp 1018054153
transform 1 0 3200 0 1 7280
box -16 -6 32 210
use FILL  FILL_459
timestamp 1018054153
transform 1 0 3216 0 1 7280
box -16 -6 32 210
use FILL  FILL_461
timestamp 1018054153
transform 1 0 3232 0 1 7280
box -16 -6 32 210
use FILL  FILL_463
timestamp 1018054153
transform 1 0 3248 0 1 7280
box -16 -6 32 210
use FILL  FILL_465
timestamp 1018054153
transform 1 0 3264 0 1 7280
box -16 -6 32 210
use FILL  FILL_467
timestamp 1018054153
transform 1 0 3280 0 1 7280
box -16 -6 32 210
use FILL  FILL_469
timestamp 1018054153
transform 1 0 3296 0 1 7280
box -16 -6 32 210
use FILL  FILL_471
timestamp 1018054153
transform 1 0 3312 0 1 7280
box -16 -6 32 210
use FILL  FILL_473
timestamp 1018054153
transform 1 0 3328 0 1 7280
box -16 -6 32 210
use FILL  FILL_475
timestamp 1018054153
transform 1 0 3344 0 1 7280
box -16 -6 32 210
use FILL  FILL_477
timestamp 1018054153
transform 1 0 3360 0 1 7280
box -16 -6 32 210
use FILL  FILL_479
timestamp 1018054153
transform 1 0 3376 0 1 7280
box -16 -6 32 210
use FILL  FILL_481
timestamp 1018054153
transform 1 0 3392 0 1 7280
box -16 -6 32 210
use FILL  FILL_483
timestamp 1018054153
transform 1 0 3408 0 1 7280
box -16 -6 32 210
use FILL  FILL_485
timestamp 1018054153
transform 1 0 3424 0 1 7280
box -16 -6 32 210
use FILL  FILL_487
timestamp 1018054153
transform 1 0 3440 0 1 7280
box -16 -6 32 210
use FILL  FILL_489
timestamp 1018054153
transform 1 0 3456 0 1 7280
box -16 -6 32 210
use FILL  FILL_491
timestamp 1018054153
transform 1 0 3472 0 1 7280
box -16 -6 32 210
use FILL  FILL_493
timestamp 1018054153
transform 1 0 3488 0 1 7280
box -16 -6 32 210
use FILL  FILL_495
timestamp 1018054153
transform 1 0 3504 0 1 7280
box -16 -6 32 210
use FILL  FILL_497
timestamp 1018054153
transform 1 0 3520 0 1 7280
box -16 -6 32 210
use FILL  FILL_499
timestamp 1018054153
transform 1 0 3536 0 1 7280
box -16 -6 32 210
use FILL  FILL_501
timestamp 1018054153
transform 1 0 3552 0 1 7280
box -16 -6 32 210
use FILL  FILL_503
timestamp 1018054153
transform 1 0 3568 0 1 7280
box -16 -6 32 210
use FILL  FILL_505
timestamp 1018054153
transform 1 0 3584 0 1 7280
box -16 -6 32 210
use FILL  FILL_507
timestamp 1018054153
transform 1 0 3600 0 1 7280
box -16 -6 32 210
use FILL  FILL_509
timestamp 1018054153
transform 1 0 3616 0 1 7280
box -16 -6 32 210
use FILL  FILL_511
timestamp 1018054153
transform 1 0 3632 0 1 7280
box -16 -6 32 210
use FILL  FILL_513
timestamp 1018054153
transform 1 0 3648 0 1 7280
box -16 -6 32 210
use FILL  FILL_515
timestamp 1018054153
transform 1 0 3664 0 1 7280
box -16 -6 32 210
use FILL  FILL_517
timestamp 1018054153
transform 1 0 3680 0 1 7280
box -16 -6 32 210
use FILL  FILL_519
timestamp 1018054153
transform 1 0 3696 0 1 7280
box -16 -6 32 210
use FILL  FILL_521
timestamp 1018054153
transform 1 0 3712 0 1 7280
box -16 -6 32 210
use FILL  FILL_523
timestamp 1018054153
transform 1 0 3728 0 1 7280
box -16 -6 32 210
use FILL  FILL_525
timestamp 1018054153
transform 1 0 3744 0 1 7280
box -16 -6 32 210
use FILL  FILL_527
timestamp 1018054153
transform 1 0 3760 0 1 7280
box -16 -6 32 210
use FILL  FILL_529
timestamp 1018054153
transform 1 0 3776 0 1 7280
box -16 -6 32 210
use FILL  FILL_531
timestamp 1018054153
transform 1 0 3792 0 1 7280
box -16 -6 32 210
use FILL  FILL_533
timestamp 1018054153
transform 1 0 3808 0 1 7280
box -16 -6 32 210
use FILL  FILL_535
timestamp 1018054153
transform 1 0 3824 0 1 7280
box -16 -6 32 210
use FILL  FILL_537
timestamp 1018054153
transform 1 0 3840 0 1 7280
box -16 -6 32 210
use FILL  FILL_539
timestamp 1018054153
transform 1 0 3856 0 1 7280
box -16 -6 32 210
use FILL  FILL_541
timestamp 1018054153
transform 1 0 3872 0 1 7280
box -16 -6 32 210
use FILL  FILL_543
timestamp 1018054153
transform 1 0 3888 0 1 7280
box -16 -6 32 210
use FILL  FILL_545
timestamp 1018054153
transform 1 0 3904 0 1 7280
box -16 -6 32 210
use FILL  FILL_547
timestamp 1018054153
transform 1 0 3920 0 1 7280
box -16 -6 32 210
use FILL  FILL_549
timestamp 1018054153
transform 1 0 3936 0 1 7280
box -16 -6 32 210
use FILL  FILL_551
timestamp 1018054153
transform 1 0 3952 0 1 7280
box -16 -6 32 210
use FILL  FILL_553
timestamp 1018054153
transform 1 0 3968 0 1 7280
box -16 -6 32 210
use FILL  FILL_555
timestamp 1018054153
transform 1 0 3984 0 1 7280
box -16 -6 32 210
use FILL  FILL_557
timestamp 1018054153
transform 1 0 4000 0 1 7280
box -16 -6 32 210
use FILL  FILL_559
timestamp 1018054153
transform 1 0 4016 0 1 7280
box -16 -6 32 210
use FILL  FILL_561
timestamp 1018054153
transform 1 0 4032 0 1 7280
box -16 -6 32 210
use FILL  FILL_563
timestamp 1018054153
transform 1 0 4048 0 1 7280
box -16 -6 32 210
use FILL  FILL_565
timestamp 1018054153
transform 1 0 4064 0 1 7280
box -16 -6 32 210
use FILL  FILL_567
timestamp 1018054153
transform 1 0 4080 0 1 7280
box -16 -6 32 210
use FILL  FILL_569
timestamp 1018054153
transform 1 0 4096 0 1 7280
box -16 -6 32 210
use FILL  FILL_571
timestamp 1018054153
transform 1 0 4112 0 1 7280
box -16 -6 32 210
use FILL  FILL_573
timestamp 1018054153
transform 1 0 4128 0 1 7280
box -16 -6 32 210
use FILL  FILL_575
timestamp 1018054153
transform 1 0 4144 0 1 7280
box -16 -6 32 210
use FILL  FILL_577
timestamp 1018054153
transform 1 0 4160 0 1 7280
box -16 -6 32 210
use FILL  FILL_579
timestamp 1018054153
transform 1 0 4176 0 1 7280
box -16 -6 32 210
use FILL  FILL_581
timestamp 1018054153
transform 1 0 4192 0 1 7280
box -16 -6 32 210
use FILL  FILL_583
timestamp 1018054153
transform 1 0 4208 0 1 7280
box -16 -6 32 210
use FILL  FILL_585
timestamp 1018054153
transform 1 0 4224 0 1 7280
box -16 -6 32 210
use FILL  FILL_587
timestamp 1018054153
transform 1 0 4240 0 1 7280
box -16 -6 32 210
use FILL  FILL_589
timestamp 1018054153
transform 1 0 4256 0 1 7280
box -16 -6 32 210
use FILL  FILL_591
timestamp 1018054153
transform 1 0 4272 0 1 7280
box -16 -6 32 210
use FILL  FILL_593
timestamp 1018054153
transform 1 0 4288 0 1 7280
box -16 -6 32 210
use FILL  FILL_595
timestamp 1018054153
transform 1 0 4304 0 1 7280
box -16 -6 32 210
use FILL  FILL_597
timestamp 1018054153
transform 1 0 4320 0 1 7280
box -16 -6 32 210
use FILL  FILL_599
timestamp 1018054153
transform 1 0 4336 0 1 7280
box -16 -6 32 210
use FILL  FILL_601
timestamp 1018054153
transform 1 0 4352 0 1 7280
box -16 -6 32 210
use FILL  FILL_603
timestamp 1018054153
transform 1 0 4368 0 1 7280
box -16 -6 32 210
use FILL  FILL_605
timestamp 1018054153
transform 1 0 4384 0 1 7280
box -16 -6 32 210
use FILL  FILL_607
timestamp 1018054153
transform 1 0 4400 0 1 7280
box -16 -6 32 210
use FILL  FILL_609
timestamp 1018054153
transform 1 0 4416 0 1 7280
box -16 -6 32 210
use FILL  FILL_611
timestamp 1018054153
transform 1 0 4432 0 1 7280
box -16 -6 32 210
use FILL  FILL_613
timestamp 1018054153
transform 1 0 4448 0 1 7280
box -16 -6 32 210
use FILL  FILL_615
timestamp 1018054153
transform 1 0 4464 0 1 7280
box -16 -6 32 210
use FILL  FILL_617
timestamp 1018054153
transform 1 0 4480 0 1 7280
box -16 -6 32 210
use FILL  FILL_619
timestamp 1018054153
transform 1 0 4496 0 1 7280
box -16 -6 32 210
use FILL  FILL_621
timestamp 1018054153
transform 1 0 4512 0 1 7280
box -16 -6 32 210
use FILL  FILL_623
timestamp 1018054153
transform 1 0 4528 0 1 7280
box -16 -6 32 210
use FILL  FILL_625
timestamp 1018054153
transform 1 0 4544 0 1 7280
box -16 -6 32 210
use FILL  FILL_627
timestamp 1018054153
transform 1 0 4560 0 1 7280
box -16 -6 32 210
use FILL  FILL_629
timestamp 1018054153
transform 1 0 4576 0 1 7280
box -16 -6 32 210
use FILL  FILL_631
timestamp 1018054153
transform 1 0 4592 0 1 7280
box -16 -6 32 210
use FILL  FILL_633
timestamp 1018054153
transform 1 0 4608 0 1 7280
box -16 -6 32 210
use FILL  FILL_635
timestamp 1018054153
transform 1 0 4624 0 1 7280
box -16 -6 32 210
use FILL  FILL_637
timestamp 1018054153
transform 1 0 4640 0 1 7280
box -16 -6 32 210
use FILL  FILL_639
timestamp 1018054153
transform 1 0 4656 0 1 7280
box -16 -6 32 210
use FILL  FILL_641
timestamp 1018054153
transform 1 0 4672 0 1 7280
box -16 -6 32 210
use FILL  FILL_643
timestamp 1018054153
transform 1 0 4688 0 1 7280
box -16 -6 32 210
use FILL  FILL_645
timestamp 1018054153
transform 1 0 4704 0 1 7280
box -16 -6 32 210
use FILL  FILL_647
timestamp 1018054153
transform 1 0 4720 0 1 7280
box -16 -6 32 210
use FILL  FILL_649
timestamp 1018054153
transform 1 0 4736 0 1 7280
box -16 -6 32 210
use FILL  FILL_651
timestamp 1018054153
transform 1 0 4752 0 1 7280
box -16 -6 32 210
use FILL  FILL_653
timestamp 1018054153
transform 1 0 4768 0 1 7280
box -16 -6 32 210
use FILL  FILL_655
timestamp 1018054153
transform 1 0 4784 0 1 7280
box -16 -6 32 210
use FILL  FILL_657
timestamp 1018054153
transform 1 0 4800 0 1 7280
box -16 -6 32 210
use FILL  FILL_659
timestamp 1018054153
transform 1 0 4816 0 1 7280
box -16 -6 32 210
use FILL  FILL_661
timestamp 1018054153
transform 1 0 4832 0 1 7280
box -16 -6 32 210
use FILL  FILL_663
timestamp 1018054153
transform 1 0 4848 0 1 7280
box -16 -6 32 210
use FILL  FILL_665
timestamp 1018054153
transform 1 0 4864 0 1 7280
box -16 -6 32 210
use FILL  FILL_667
timestamp 1018054153
transform 1 0 4880 0 1 7280
box -16 -6 32 210
use FILL  FILL_669
timestamp 1018054153
transform 1 0 4896 0 1 7280
box -16 -6 32 210
use FILL  FILL_671
timestamp 1018054153
transform 1 0 4912 0 1 7280
box -16 -6 32 210
use FILL  FILL_673
timestamp 1018054153
transform 1 0 4928 0 1 7280
box -16 -6 32 210
use FILL  FILL_675
timestamp 1018054153
transform 1 0 4944 0 1 7280
box -16 -6 32 210
use FILL  FILL_677
timestamp 1018054153
transform 1 0 4960 0 1 7280
box -16 -6 32 210
use FILL  FILL_679
timestamp 1018054153
transform 1 0 4976 0 1 7280
box -16 -6 32 210
use FILL  FILL_681
timestamp 1018054153
transform 1 0 4992 0 1 7280
box -16 -6 32 210
use FILL  FILL_683
timestamp 1018054153
transform 1 0 5008 0 1 7280
box -16 -6 32 210
use FILL  FILL_685
timestamp 1018054153
transform 1 0 5024 0 1 7280
box -16 -6 32 210
use FILL  FILL_687
timestamp 1018054153
transform 1 0 5040 0 1 7280
box -16 -6 32 210
use FILL  FILL_689
timestamp 1018054153
transform 1 0 5056 0 1 7280
box -16 -6 32 210
use FILL  FILL_691
timestamp 1018054153
transform 1 0 5072 0 1 7280
box -16 -6 32 210
use FILL  FILL_693
timestamp 1018054153
transform 1 0 5088 0 1 7280
box -16 -6 32 210
use FILL  FILL_695
timestamp 1018054153
transform 1 0 5104 0 1 7280
box -16 -6 32 210
use FILL  FILL_697
timestamp 1018054153
transform 1 0 5120 0 1 7280
box -16 -6 32 210
use FILL  FILL_699
timestamp 1018054153
transform 1 0 5136 0 1 7280
box -16 -6 32 210
use FILL  FILL_701
timestamp 1018054153
transform 1 0 5152 0 1 7280
box -16 -6 32 210
use FILL  FILL_703
timestamp 1018054153
transform 1 0 5168 0 1 7280
box -16 -6 32 210
use FILL  FILL_705
timestamp 1018054153
transform 1 0 5184 0 1 7280
box -16 -6 32 210
use FILL  FILL_707
timestamp 1018054153
transform 1 0 5200 0 1 7280
box -16 -6 32 210
use FILL  FILL_709
timestamp 1018054153
transform 1 0 5216 0 1 7280
box -16 -6 32 210
use FILL  FILL_711
timestamp 1018054153
transform 1 0 5232 0 1 7280
box -16 -6 32 210
use FILL  FILL_713
timestamp 1018054153
transform 1 0 5248 0 1 7280
box -16 -6 32 210
use FILL  FILL_715
timestamp 1018054153
transform 1 0 5264 0 1 7280
box -16 -6 32 210
use FILL  FILL_717
timestamp 1018054153
transform 1 0 5280 0 1 7280
box -16 -6 32 210
use FILL  FILL_719
timestamp 1018054153
transform 1 0 5296 0 1 7280
box -16 -6 32 210
use FILL  FILL_721
timestamp 1018054153
transform 1 0 5312 0 1 7280
box -16 -6 32 210
use FILL  FILL_723
timestamp 1018054153
transform 1 0 5328 0 1 7280
box -16 -6 32 210
use FILL  FILL_725
timestamp 1018054153
transform 1 0 5344 0 1 7280
box -16 -6 32 210
use FILL  FILL_727
timestamp 1018054153
transform 1 0 5360 0 1 7280
box -16 -6 32 210
use FILL  FILL_729
timestamp 1018054153
transform 1 0 5376 0 1 7280
box -16 -6 32 210
use FILL  FILL_731
timestamp 1018054153
transform 1 0 5392 0 1 7280
box -16 -6 32 210
use FILL  FILL_733
timestamp 1018054153
transform 1 0 5408 0 1 7280
box -16 -6 32 210
use FILL  FILL_735
timestamp 1018054153
transform 1 0 5424 0 1 7280
box -16 -6 32 210
use FILL  FILL_737
timestamp 1018054153
transform 1 0 5440 0 1 7280
box -16 -6 32 210
use FILL  FILL_739
timestamp 1018054153
transform 1 0 5456 0 1 7280
box -16 -6 32 210
use FILL  FILL_741
timestamp 1018054153
transform 1 0 5472 0 1 7280
box -16 -6 32 210
use FILL  FILL_743
timestamp 1018054153
transform 1 0 5488 0 1 7280
box -16 -6 32 210
use FILL  FILL_745
timestamp 1018054153
transform 1 0 5504 0 1 7280
box -16 -6 32 210
use FILL  FILL_747
timestamp 1018054153
transform 1 0 5520 0 1 7280
box -16 -6 32 210
use FILL  FILL_749
timestamp 1018054153
transform 1 0 5536 0 1 7280
box -16 -6 32 210
use FILL  FILL_751
timestamp 1018054153
transform 1 0 5552 0 1 7280
box -16 -6 32 210
use FILL  FILL_753
timestamp 1018054153
transform 1 0 5568 0 1 7280
box -16 -6 32 210
use FILL  FILL_755
timestamp 1018054153
transform 1 0 5584 0 1 7280
box -16 -6 32 210
use FILL  FILL_757
timestamp 1018054153
transform 1 0 5600 0 1 7280
box -16 -6 32 210
use FILL  FILL_759
timestamp 1018054153
transform 1 0 5616 0 1 7280
box -16 -6 32 210
use FILL  FILL_761
timestamp 1018054153
transform 1 0 5632 0 1 7280
box -16 -6 32 210
use FILL  FILL_763
timestamp 1018054153
transform 1 0 5648 0 1 7280
box -16 -6 32 210
use FILL  FILL_765
timestamp 1018054153
transform 1 0 5664 0 1 7280
box -16 -6 32 210
use FILL  FILL_767
timestamp 1018054153
transform 1 0 5680 0 1 7280
box -16 -6 32 210
use FILL  FILL_769
timestamp 1018054153
transform 1 0 5696 0 1 7280
box -16 -6 32 210
use FILL  FILL_771
timestamp 1018054153
transform 1 0 5712 0 1 7280
box -16 -6 32 210
use FILL  FILL_773
timestamp 1018054153
transform 1 0 5728 0 1 7280
box -16 -6 32 210
use FILL  FILL_775
timestamp 1018054153
transform 1 0 5744 0 1 7280
box -16 -6 32 210
use FILL  FILL_777
timestamp 1018054153
transform 1 0 5760 0 1 7280
box -16 -6 32 210
use FILL  FILL_779
timestamp 1018054153
transform 1 0 5776 0 1 7280
box -16 -6 32 210
use FILL  FILL_781
timestamp 1018054153
transform 1 0 5792 0 1 7280
box -16 -6 32 210
use FILL  FILL_783
timestamp 1018054153
transform 1 0 5808 0 1 7280
box -16 -6 32 210
use FILL  FILL_785
timestamp 1018054153
transform 1 0 5824 0 1 7280
box -16 -6 32 210
use FILL  FILL_787
timestamp 1018054153
transform 1 0 5840 0 1 7280
box -16 -6 32 210
use FILL  FILL_789
timestamp 1018054153
transform 1 0 5856 0 1 7280
box -16 -6 32 210
use FILL  FILL_791
timestamp 1018054153
transform 1 0 5872 0 1 7280
box -16 -6 32 210
use FILL  FILL_793
timestamp 1018054153
transform 1 0 5888 0 1 7280
box -16 -6 32 210
use FILL  FILL_795
timestamp 1018054153
transform 1 0 5904 0 1 7280
box -16 -6 32 210
use FILL  FILL_797
timestamp 1018054153
transform 1 0 5920 0 1 7280
box -16 -6 32 210
use FILL  FILL_799
timestamp 1018054153
transform 1 0 5936 0 1 7280
box -16 -6 32 210
use FILL  FILL_801
timestamp 1018054153
transform 1 0 5952 0 1 7280
box -16 -6 32 210
use FILL  FILL_803
timestamp 1018054153
transform 1 0 5968 0 1 7280
box -16 -6 32 210
use FILL  FILL_805
timestamp 1018054153
transform 1 0 5984 0 1 7280
box -16 -6 32 210
use FILL  FILL_807
timestamp 1018054153
transform 1 0 6000 0 1 7280
box -16 -6 32 210
use FILL  FILL_809
timestamp 1018054153
transform 1 0 6016 0 1 7280
box -16 -6 32 210
use FILL  FILL_811
timestamp 1018054153
transform 1 0 6032 0 1 7280
box -16 -6 32 210
use FILL  FILL_813
timestamp 1018054153
transform 1 0 6048 0 1 7280
box -16 -6 32 210
use FILL  FILL_815
timestamp 1018054153
transform 1 0 6064 0 1 7280
box -16 -6 32 210
use FILL  FILL_817
timestamp 1018054153
transform 1 0 6080 0 1 7280
box -16 -6 32 210
use FILL  FILL_819
timestamp 1018054153
transform 1 0 6096 0 1 7280
box -16 -6 32 210
use FILL  FILL_821
timestamp 1018054153
transform 1 0 6112 0 1 7280
box -16 -6 32 210
use FILL  FILL_823
timestamp 1018054153
transform 1 0 6128 0 1 7280
box -16 -6 32 210
use FILL  FILL_825
timestamp 1018054153
transform 1 0 6144 0 1 7280
box -16 -6 32 210
use FILL  FILL_827
timestamp 1018054153
transform 1 0 6160 0 1 7280
box -16 -6 32 210
use FILL  FILL_829
timestamp 1018054153
transform 1 0 6176 0 1 7280
box -16 -6 32 210
use FILL  FILL_831
timestamp 1018054153
transform 1 0 6192 0 1 7280
box -16 -6 32 210
use FILL  FILL_833
timestamp 1018054153
transform 1 0 6208 0 1 7280
box -16 -6 32 210
use FILL  FILL_835
timestamp 1018054153
transform 1 0 6224 0 1 7280
box -16 -6 32 210
use FILL  FILL_837
timestamp 1018054153
transform 1 0 6240 0 1 7280
box -16 -6 32 210
use FILL  FILL_839
timestamp 1018054153
transform 1 0 6256 0 1 7280
box -16 -6 32 210
use FILL  FILL_841
timestamp 1018054153
transform 1 0 6272 0 1 7280
box -16 -6 32 210
use FILL  FILL_843
timestamp 1018054153
transform 1 0 6288 0 1 7280
box -16 -6 32 210
use FILL  FILL_845
timestamp 1018054153
transform 1 0 6304 0 1 7280
box -16 -6 32 210
use FILL  FILL_847
timestamp 1018054153
transform 1 0 6320 0 1 7280
box -16 -6 32 210
use FILL  FILL_849
timestamp 1018054153
transform 1 0 6336 0 1 7280
box -16 -6 32 210
use FILL  FILL_851
timestamp 1018054153
transform 1 0 6352 0 1 7280
box -16 -6 32 210
use FILL  FILL_853
timestamp 1018054153
transform 1 0 6368 0 1 7280
box -16 -6 32 210
use FILL  FILL_855
timestamp 1018054153
transform 1 0 6384 0 1 7280
box -16 -6 32 210
use FILL  FILL_857
timestamp 1018054153
transform 1 0 6400 0 1 7280
box -16 -6 32 210
use FILL  FILL_859
timestamp 1018054153
transform 1 0 6416 0 1 7280
box -16 -6 32 210
use FILL  FILL_861
timestamp 1018054153
transform 1 0 6432 0 1 7280
box -16 -6 32 210
use FILL  FILL_863
timestamp 1018054153
transform 1 0 6448 0 1 7280
box -16 -6 32 210
use FILL  FILL_865
timestamp 1018054153
transform 1 0 6464 0 1 7280
box -16 -6 32 210
use FILL  FILL_867
timestamp 1018054153
transform 1 0 6480 0 1 7280
box -16 -6 32 210
use FILL  FILL_869
timestamp 1018054153
transform 1 0 6496 0 1 7280
box -16 -6 32 210
use FILL  FILL_871
timestamp 1018054153
transform 1 0 6512 0 1 7280
box -16 -6 32 210
use FILL  FILL_873
timestamp 1018054153
transform 1 0 6528 0 1 7280
box -16 -6 32 210
use FILL  FILL_875
timestamp 1018054153
transform 1 0 6544 0 1 7280
box -16 -6 32 210
use FILL  FILL_877
timestamp 1018054153
transform 1 0 6560 0 1 7280
box -16 -6 32 210
use FILL  FILL_879
timestamp 1018054153
transform 1 0 6576 0 1 7280
box -16 -6 32 210
use FILL  FILL_881
timestamp 1018054153
transform 1 0 6592 0 1 7280
box -16 -6 32 210
use FILL  FILL_883
timestamp 1018054153
transform 1 0 6608 0 1 7280
box -16 -6 32 210
use FILL  FILL_885
timestamp 1018054153
transform 1 0 6624 0 1 7280
box -16 -6 32 210
use FILL  FILL_887
timestamp 1018054153
transform 1 0 6640 0 1 7280
box -16 -6 32 210
use FILL  FILL_889
timestamp 1018054153
transform 1 0 6656 0 1 7280
box -16 -6 32 210
use FILL  FILL_891
timestamp 1018054153
transform 1 0 6672 0 1 7280
box -16 -6 32 210
use FILL  FILL_893
timestamp 1018054153
transform 1 0 6688 0 1 7280
box -16 -6 32 210
use FILL  FILL_895
timestamp 1018054153
transform 1 0 6704 0 1 7280
box -16 -6 32 210
use FILL  FILL_897
timestamp 1018054153
transform 1 0 6720 0 1 7280
box -16 -6 32 210
use FILL  FILL_899
timestamp 1018054153
transform 1 0 6736 0 1 7280
box -16 -6 32 210
use FILL  FILL_901
timestamp 1018054153
transform 1 0 6752 0 1 7280
box -16 -6 32 210
use FILL  FILL_903
timestamp 1018054153
transform 1 0 6768 0 1 7280
box -16 -6 32 210
use FILL  FILL_905
timestamp 1018054153
transform 1 0 6784 0 1 7280
box -16 -6 32 210
use FILL  FILL_907
timestamp 1018054153
transform 1 0 6800 0 1 7280
box -16 -6 32 210
use FILL  FILL_909
timestamp 1018054153
transform 1 0 6816 0 1 7280
box -16 -6 32 210
use FILL  FILL_911
timestamp 1018054153
transform 1 0 6832 0 1 7280
box -16 -6 32 210
use FILL  FILL_913
timestamp 1018054153
transform 1 0 6848 0 1 7280
box -16 -6 32 210
use FILL  FILL_915
timestamp 1018054153
transform 1 0 6864 0 1 7280
box -16 -6 32 210
use FILL  FILL_917
timestamp 1018054153
transform 1 0 6880 0 1 7280
box -16 -6 32 210
use FILL  FILL_919
timestamp 1018054153
transform 1 0 6896 0 1 7280
box -16 -6 32 210
use FILL  FILL_921
timestamp 1018054153
transform 1 0 6912 0 1 7280
box -16 -6 32 210
use FILL  FILL_923
timestamp 1018054153
transform 1 0 6928 0 1 7280
box -16 -6 32 210
use FILL  FILL_925
timestamp 1018054153
transform 1 0 6944 0 1 7280
box -16 -6 32 210
use FILL  FILL_927
timestamp 1018054153
transform 1 0 6960 0 1 7280
box -16 -6 32 210
use FILL  FILL_929
timestamp 1018054153
transform 1 0 6976 0 1 7280
box -16 -6 32 210
use FILL  FILL_931
timestamp 1018054153
transform 1 0 6992 0 1 7280
box -16 -6 32 210
use FILL  FILL_933
timestamp 1018054153
transform 1 0 7008 0 1 7280
box -16 -6 32 210
use FILL  FILL_935
timestamp 1018054153
transform 1 0 7024 0 1 7280
box -16 -6 32 210
use FILL  FILL_937
timestamp 1018054153
transform 1 0 7040 0 1 7280
box -16 -6 32 210
use FILL  FILL_939
timestamp 1018054153
transform 1 0 7056 0 1 7280
box -16 -6 32 210
use FILL  FILL_941
timestamp 1018054153
transform 1 0 7072 0 1 7280
box -16 -6 32 210
use FILL  FILL_943
timestamp 1018054153
transform 1 0 7088 0 1 7280
box -16 -6 32 210
use FILL  FILL_945
timestamp 1018054153
transform 1 0 7104 0 1 7280
box -16 -6 32 210
use FILL  FILL_947
timestamp 1018054153
transform 1 0 7120 0 1 7280
box -16 -6 32 210
use FILL  FILL_949
timestamp 1018054153
transform 1 0 7136 0 1 7280
box -16 -6 32 210
use FILL  FILL_951
timestamp 1018054153
transform 1 0 7152 0 1 7280
box -16 -6 32 210
use FILL  FILL_953
timestamp 1018054153
transform 1 0 7168 0 1 7280
box -16 -6 32 210
use FILL  FILL_955
timestamp 1018054153
transform 1 0 7184 0 1 7280
box -16 -6 32 210
use FILL  FILL_957
timestamp 1018054153
transform 1 0 7200 0 1 7280
box -16 -6 32 210
use FILL  FILL_959
timestamp 1018054153
transform 1 0 7216 0 1 7280
box -16 -6 32 210
use FILL  FILL_961
timestamp 1018054153
transform 1 0 7232 0 1 7280
box -16 -6 32 210
use FILL  FILL_963
timestamp 1018054153
transform 1 0 7248 0 1 7280
box -16 -6 32 210
use FILL  FILL_965
timestamp 1018054153
transform 1 0 7264 0 1 7280
box -16 -6 32 210
use FILL  FILL_967
timestamp 1018054153
transform 1 0 7280 0 1 7280
box -16 -6 32 210
use FILL  FILL_969
timestamp 1018054153
transform 1 0 7296 0 1 7280
box -16 -6 32 210
use FILL  FILL_971
timestamp 1018054153
transform 1 0 7312 0 1 7280
box -16 -6 32 210
use FILL  FILL_973
timestamp 1018054153
transform 1 0 7328 0 1 7280
box -16 -6 32 210
use FILL  FILL_975
timestamp 1018054153
transform 1 0 7344 0 1 7280
box -16 -6 32 210
use FILL  FILL_977
timestamp 1018054153
transform 1 0 7360 0 1 7280
box -16 -6 32 210
use FILL  FILL_979
timestamp 1018054153
transform 1 0 7376 0 1 7280
box -16 -6 32 210
use FILL  FILL_981
timestamp 1018054153
transform 1 0 7392 0 1 7280
box -16 -6 32 210
use FILL  FILL_983
timestamp 1018054153
transform 1 0 7408 0 1 7280
box -16 -6 32 210
use FILL  FILL_985
timestamp 1018054153
transform 1 0 7424 0 1 7280
box -16 -6 32 210
use FILL  FILL_987
timestamp 1018054153
transform 1 0 7440 0 1 7280
box -16 -6 32 210
use FILL  FILL_989
timestamp 1018054153
transform 1 0 7456 0 1 7280
box -16 -6 32 210
use FILL  FILL_991
timestamp 1018054153
transform 1 0 7472 0 1 7280
box -16 -6 32 210
use FILL  FILL_993
timestamp 1018054153
transform 1 0 7488 0 1 7280
box -16 -6 32 210
use FILL  FILL_995
timestamp 1018054153
transform 1 0 7504 0 1 7280
box -16 -6 32 210
use FILL  FILL_997
timestamp 1018054153
transform 1 0 7520 0 1 7280
box -16 -6 32 210
use FILL  FILL_999
timestamp 1018054153
transform 1 0 7536 0 1 7280
box -16 -6 32 210
use FILL  FILL_1001
timestamp 1018054153
transform 1 0 7552 0 1 7280
box -16 -6 32 210
use FILL  FILL_1003
timestamp 1018054153
transform 1 0 7568 0 1 7280
box -16 -6 32 210
use FILL  FILL_1005
timestamp 1018054153
transform 1 0 7584 0 1 7280
box -16 -6 32 210
use FILL  FILL_1007
timestamp 1018054153
transform 1 0 7600 0 1 7280
box -16 -6 32 210
use FILL  FILL_1009
timestamp 1018054153
transform 1 0 7616 0 1 7280
box -16 -6 32 210
use FILL  FILL_1011
timestamp 1018054153
transform 1 0 7632 0 1 7280
box -16 -6 32 210
use FILL  FILL_1013
timestamp 1018054153
transform 1 0 7648 0 1 7280
box -16 -6 32 210
use FILL  FILL_1015
timestamp 1018054153
transform 1 0 7664 0 1 7280
box -16 -6 32 210
use FILL  FILL_1017
timestamp 1018054153
transform 1 0 7680 0 1 7280
box -16 -6 32 210
use FILL  FILL_1019
timestamp 1018054153
transform 1 0 7696 0 1 7280
box -16 -6 32 210
use FILL  FILL_1021
timestamp 1018054153
transform 1 0 7712 0 1 7280
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_3
timestamp 1542725905
transform 1 0 7908 0 1 7280
box -48 -6 48 6
use FILL  FILL_342
timestamp 1018054153
transform 1 0 2272 0 -1 7280
box -16 -6 32 210
use FILL  FILL_344
timestamp 1018054153
transform 1 0 2288 0 -1 7280
box -16 -6 32 210
use FILL  FILL_346
timestamp 1018054153
transform 1 0 2304 0 -1 7280
box -16 -6 32 210
use FILL  FILL_348
timestamp 1018054153
transform 1 0 2320 0 -1 7280
box -16 -6 32 210
use FILL  FILL_350
timestamp 1018054153
transform 1 0 2336 0 -1 7280
box -16 -6 32 210
use FILL  FILL_352
timestamp 1018054153
transform 1 0 2352 0 -1 7280
box -16 -6 32 210
use FILL  FILL_354
timestamp 1018054153
transform 1 0 2368 0 -1 7280
box -16 -6 32 210
use FILL  FILL_356
timestamp 1018054153
transform 1 0 2384 0 -1 7280
box -16 -6 32 210
use FILL  FILL_358
timestamp 1018054153
transform 1 0 2400 0 -1 7280
box -16 -6 32 210
use FILL  FILL_360
timestamp 1018054153
transform 1 0 2416 0 -1 7280
box -16 -6 32 210
use FILL  FILL_362
timestamp 1018054153
transform 1 0 2432 0 -1 7280
box -16 -6 32 210
use FILL  FILL_364
timestamp 1018054153
transform 1 0 2448 0 -1 7280
box -16 -6 32 210
use FILL  FILL_366
timestamp 1018054153
transform 1 0 2464 0 -1 7280
box -16 -6 32 210
use FILL  FILL_368
timestamp 1018054153
transform 1 0 2480 0 -1 7280
box -16 -6 32 210
use FILL  FILL_370
timestamp 1018054153
transform 1 0 2496 0 -1 7280
box -16 -6 32 210
use FILL  FILL_372
timestamp 1018054153
transform 1 0 2512 0 -1 7280
box -16 -6 32 210
use FILL  FILL_374
timestamp 1018054153
transform 1 0 2528 0 -1 7280
box -16 -6 32 210
use FILL  FILL_376
timestamp 1018054153
transform 1 0 2544 0 -1 7280
box -16 -6 32 210
use FILL  FILL_378
timestamp 1018054153
transform 1 0 2560 0 -1 7280
box -16 -6 32 210
use FILL  FILL_380
timestamp 1018054153
transform 1 0 2576 0 -1 7280
box -16 -6 32 210
use FILL  FILL_382
timestamp 1018054153
transform 1 0 2592 0 -1 7280
box -16 -6 32 210
use FILL  FILL_384
timestamp 1018054153
transform 1 0 2608 0 -1 7280
box -16 -6 32 210
use FILL  FILL_386
timestamp 1018054153
transform 1 0 2624 0 -1 7280
box -16 -6 32 210
use FILL  FILL_388
timestamp 1018054153
transform 1 0 2640 0 -1 7280
box -16 -6 32 210
use FILL  FILL_390
timestamp 1018054153
transform 1 0 2656 0 -1 7280
box -16 -6 32 210
use FILL  FILL_392
timestamp 1018054153
transform 1 0 2672 0 -1 7280
box -16 -6 32 210
use FILL  FILL_394
timestamp 1018054153
transform 1 0 2688 0 -1 7280
box -16 -6 32 210
use FILL  FILL_396
timestamp 1018054153
transform 1 0 2704 0 -1 7280
box -16 -6 32 210
use FILL  FILL_398
timestamp 1018054153
transform 1 0 2720 0 -1 7280
box -16 -6 32 210
use FILL  FILL_400
timestamp 1018054153
transform 1 0 2736 0 -1 7280
box -16 -6 32 210
use FILL  FILL_402
timestamp 1018054153
transform 1 0 2752 0 -1 7280
box -16 -6 32 210
use FILL  FILL_404
timestamp 1018054153
transform 1 0 2768 0 -1 7280
box -16 -6 32 210
use FILL  FILL_406
timestamp 1018054153
transform 1 0 2784 0 -1 7280
box -16 -6 32 210
use FILL  FILL_408
timestamp 1018054153
transform 1 0 2800 0 -1 7280
box -16 -6 32 210
use FILL  FILL_410
timestamp 1018054153
transform 1 0 2816 0 -1 7280
box -16 -6 32 210
use FILL  FILL_412
timestamp 1018054153
transform 1 0 2832 0 -1 7280
box -16 -6 32 210
use FILL  FILL_414
timestamp 1018054153
transform 1 0 2848 0 -1 7280
box -16 -6 32 210
use FILL  FILL_416
timestamp 1018054153
transform 1 0 2864 0 -1 7280
box -16 -6 32 210
use FILL  FILL_418
timestamp 1018054153
transform 1 0 2880 0 -1 7280
box -16 -6 32 210
use FILL  FILL_420
timestamp 1018054153
transform 1 0 2896 0 -1 7280
box -16 -6 32 210
use FILL  FILL_422
timestamp 1018054153
transform 1 0 2912 0 -1 7280
box -16 -6 32 210
use FILL  FILL_424
timestamp 1018054153
transform 1 0 2928 0 -1 7280
box -16 -6 32 210
use FILL  FILL_426
timestamp 1018054153
transform 1 0 2944 0 -1 7280
box -16 -6 32 210
use FILL  FILL_428
timestamp 1018054153
transform 1 0 2960 0 -1 7280
box -16 -6 32 210
use FILL  FILL_430
timestamp 1018054153
transform 1 0 2976 0 -1 7280
box -16 -6 32 210
use FILL  FILL_432
timestamp 1018054153
transform 1 0 2992 0 -1 7280
box -16 -6 32 210
use FILL  FILL_434
timestamp 1018054153
transform 1 0 3008 0 -1 7280
box -16 -6 32 210
use FILL  FILL_436
timestamp 1018054153
transform 1 0 3024 0 -1 7280
box -16 -6 32 210
use FILL  FILL_438
timestamp 1018054153
transform 1 0 3040 0 -1 7280
box -16 -6 32 210
use FILL  FILL_440
timestamp 1018054153
transform 1 0 3056 0 -1 7280
box -16 -6 32 210
use FILL  FILL_442
timestamp 1018054153
transform 1 0 3072 0 -1 7280
box -16 -6 32 210
use FILL  FILL_444
timestamp 1018054153
transform 1 0 3088 0 -1 7280
box -16 -6 32 210
use FILL  FILL_446
timestamp 1018054153
transform 1 0 3104 0 -1 7280
box -16 -6 32 210
use FILL  FILL_448
timestamp 1018054153
transform 1 0 3120 0 -1 7280
box -16 -6 32 210
use FILL  FILL_450
timestamp 1018054153
transform 1 0 3136 0 -1 7280
box -16 -6 32 210
use FILL  FILL_452
timestamp 1018054153
transform 1 0 3152 0 -1 7280
box -16 -6 32 210
use FILL  FILL_454
timestamp 1018054153
transform 1 0 3168 0 -1 7280
box -16 -6 32 210
use FILL  FILL_456
timestamp 1018054153
transform 1 0 3184 0 -1 7280
box -16 -6 32 210
use FILL  FILL_458
timestamp 1018054153
transform 1 0 3200 0 -1 7280
box -16 -6 32 210
use FILL  FILL_460
timestamp 1018054153
transform 1 0 3216 0 -1 7280
box -16 -6 32 210
use FILL  FILL_462
timestamp 1018054153
transform 1 0 3232 0 -1 7280
box -16 -6 32 210
use FILL  FILL_464
timestamp 1018054153
transform 1 0 3248 0 -1 7280
box -16 -6 32 210
use FILL  FILL_466
timestamp 1018054153
transform 1 0 3264 0 -1 7280
box -16 -6 32 210
use FILL  FILL_468
timestamp 1018054153
transform 1 0 3280 0 -1 7280
box -16 -6 32 210
use FILL  FILL_470
timestamp 1018054153
transform 1 0 3296 0 -1 7280
box -16 -6 32 210
use FILL  FILL_472
timestamp 1018054153
transform 1 0 3312 0 -1 7280
box -16 -6 32 210
use FILL  FILL_474
timestamp 1018054153
transform 1 0 3328 0 -1 7280
box -16 -6 32 210
use FILL  FILL_476
timestamp 1018054153
transform 1 0 3344 0 -1 7280
box -16 -6 32 210
use FILL  FILL_478
timestamp 1018054153
transform 1 0 3360 0 -1 7280
box -16 -6 32 210
use FILL  FILL_480
timestamp 1018054153
transform 1 0 3376 0 -1 7280
box -16 -6 32 210
use FILL  FILL_482
timestamp 1018054153
transform 1 0 3392 0 -1 7280
box -16 -6 32 210
use FILL  FILL_484
timestamp 1018054153
transform 1 0 3408 0 -1 7280
box -16 -6 32 210
use FILL  FILL_486
timestamp 1018054153
transform 1 0 3424 0 -1 7280
box -16 -6 32 210
use FILL  FILL_488
timestamp 1018054153
transform 1 0 3440 0 -1 7280
box -16 -6 32 210
use FILL  FILL_490
timestamp 1018054153
transform 1 0 3456 0 -1 7280
box -16 -6 32 210
use FILL  FILL_492
timestamp 1018054153
transform 1 0 3472 0 -1 7280
box -16 -6 32 210
use FILL  FILL_494
timestamp 1018054153
transform 1 0 3488 0 -1 7280
box -16 -6 32 210
use FILL  FILL_496
timestamp 1018054153
transform 1 0 3504 0 -1 7280
box -16 -6 32 210
use FILL  FILL_498
timestamp 1018054153
transform 1 0 3520 0 -1 7280
box -16 -6 32 210
use FILL  FILL_500
timestamp 1018054153
transform 1 0 3536 0 -1 7280
box -16 -6 32 210
use FILL  FILL_502
timestamp 1018054153
transform 1 0 3552 0 -1 7280
box -16 -6 32 210
use FILL  FILL_504
timestamp 1018054153
transform 1 0 3568 0 -1 7280
box -16 -6 32 210
use FILL  FILL_506
timestamp 1018054153
transform 1 0 3584 0 -1 7280
box -16 -6 32 210
use FILL  FILL_508
timestamp 1018054153
transform 1 0 3600 0 -1 7280
box -16 -6 32 210
use FILL  FILL_510
timestamp 1018054153
transform 1 0 3616 0 -1 7280
box -16 -6 32 210
use FILL  FILL_512
timestamp 1018054153
transform 1 0 3632 0 -1 7280
box -16 -6 32 210
use FILL  FILL_514
timestamp 1018054153
transform 1 0 3648 0 -1 7280
box -16 -6 32 210
use FILL  FILL_516
timestamp 1018054153
transform 1 0 3664 0 -1 7280
box -16 -6 32 210
use FILL  FILL_518
timestamp 1018054153
transform 1 0 3680 0 -1 7280
box -16 -6 32 210
use FILL  FILL_520
timestamp 1018054153
transform 1 0 3696 0 -1 7280
box -16 -6 32 210
use FILL  FILL_522
timestamp 1018054153
transform 1 0 3712 0 -1 7280
box -16 -6 32 210
use FILL  FILL_524
timestamp 1018054153
transform 1 0 3728 0 -1 7280
box -16 -6 32 210
use FILL  FILL_526
timestamp 1018054153
transform 1 0 3744 0 -1 7280
box -16 -6 32 210
use FILL  FILL_528
timestamp 1018054153
transform 1 0 3760 0 -1 7280
box -16 -6 32 210
use FILL  FILL_530
timestamp 1018054153
transform 1 0 3776 0 -1 7280
box -16 -6 32 210
use FILL  FILL_532
timestamp 1018054153
transform 1 0 3792 0 -1 7280
box -16 -6 32 210
use FILL  FILL_534
timestamp 1018054153
transform 1 0 3808 0 -1 7280
box -16 -6 32 210
use FILL  FILL_536
timestamp 1018054153
transform 1 0 3824 0 -1 7280
box -16 -6 32 210
use FILL  FILL_538
timestamp 1018054153
transform 1 0 3840 0 -1 7280
box -16 -6 32 210
use FILL  FILL_540
timestamp 1018054153
transform 1 0 3856 0 -1 7280
box -16 -6 32 210
use FILL  FILL_542
timestamp 1018054153
transform 1 0 3872 0 -1 7280
box -16 -6 32 210
use FILL  FILL_544
timestamp 1018054153
transform 1 0 3888 0 -1 7280
box -16 -6 32 210
use FILL  FILL_546
timestamp 1018054153
transform 1 0 3904 0 -1 7280
box -16 -6 32 210
use FILL  FILL_548
timestamp 1018054153
transform 1 0 3920 0 -1 7280
box -16 -6 32 210
use FILL  FILL_550
timestamp 1018054153
transform 1 0 3936 0 -1 7280
box -16 -6 32 210
use FILL  FILL_552
timestamp 1018054153
transform 1 0 3952 0 -1 7280
box -16 -6 32 210
use FILL  FILL_554
timestamp 1018054153
transform 1 0 3968 0 -1 7280
box -16 -6 32 210
use FILL  FILL_556
timestamp 1018054153
transform 1 0 3984 0 -1 7280
box -16 -6 32 210
use FILL  FILL_558
timestamp 1018054153
transform 1 0 4000 0 -1 7280
box -16 -6 32 210
use FILL  FILL_560
timestamp 1018054153
transform 1 0 4016 0 -1 7280
box -16 -6 32 210
use FILL  FILL_562
timestamp 1018054153
transform 1 0 4032 0 -1 7280
box -16 -6 32 210
use FILL  FILL_564
timestamp 1018054153
transform 1 0 4048 0 -1 7280
box -16 -6 32 210
use FILL  FILL_566
timestamp 1018054153
transform 1 0 4064 0 -1 7280
box -16 -6 32 210
use FILL  FILL_568
timestamp 1018054153
transform 1 0 4080 0 -1 7280
box -16 -6 32 210
use FILL  FILL_570
timestamp 1018054153
transform 1 0 4096 0 -1 7280
box -16 -6 32 210
use FILL  FILL_572
timestamp 1018054153
transform 1 0 4112 0 -1 7280
box -16 -6 32 210
use FILL  FILL_574
timestamp 1018054153
transform 1 0 4128 0 -1 7280
box -16 -6 32 210
use FILL  FILL_576
timestamp 1018054153
transform 1 0 4144 0 -1 7280
box -16 -6 32 210
use FILL  FILL_578
timestamp 1018054153
transform 1 0 4160 0 -1 7280
box -16 -6 32 210
use FILL  FILL_580
timestamp 1018054153
transform 1 0 4176 0 -1 7280
box -16 -6 32 210
use FILL  FILL_582
timestamp 1018054153
transform 1 0 4192 0 -1 7280
box -16 -6 32 210
use FILL  FILL_584
timestamp 1018054153
transform 1 0 4208 0 -1 7280
box -16 -6 32 210
use FILL  FILL_586
timestamp 1018054153
transform 1 0 4224 0 -1 7280
box -16 -6 32 210
use FILL  FILL_588
timestamp 1018054153
transform 1 0 4240 0 -1 7280
box -16 -6 32 210
use FILL  FILL_590
timestamp 1018054153
transform 1 0 4256 0 -1 7280
box -16 -6 32 210
use FILL  FILL_592
timestamp 1018054153
transform 1 0 4272 0 -1 7280
box -16 -6 32 210
use FILL  FILL_594
timestamp 1018054153
transform 1 0 4288 0 -1 7280
box -16 -6 32 210
use FILL  FILL_596
timestamp 1018054153
transform 1 0 4304 0 -1 7280
box -16 -6 32 210
use FILL  FILL_598
timestamp 1018054153
transform 1 0 4320 0 -1 7280
box -16 -6 32 210
use FILL  FILL_600
timestamp 1018054153
transform 1 0 4336 0 -1 7280
box -16 -6 32 210
use FILL  FILL_602
timestamp 1018054153
transform 1 0 4352 0 -1 7280
box -16 -6 32 210
use FILL  FILL_604
timestamp 1018054153
transform 1 0 4368 0 -1 7280
box -16 -6 32 210
use FILL  FILL_606
timestamp 1018054153
transform 1 0 4384 0 -1 7280
box -16 -6 32 210
use FILL  FILL_608
timestamp 1018054153
transform 1 0 4400 0 -1 7280
box -16 -6 32 210
use FILL  FILL_610
timestamp 1018054153
transform 1 0 4416 0 -1 7280
box -16 -6 32 210
use FILL  FILL_612
timestamp 1018054153
transform 1 0 4432 0 -1 7280
box -16 -6 32 210
use FILL  FILL_614
timestamp 1018054153
transform 1 0 4448 0 -1 7280
box -16 -6 32 210
use FILL  FILL_616
timestamp 1018054153
transform 1 0 4464 0 -1 7280
box -16 -6 32 210
use FILL  FILL_618
timestamp 1018054153
transform 1 0 4480 0 -1 7280
box -16 -6 32 210
use FILL  FILL_620
timestamp 1018054153
transform 1 0 4496 0 -1 7280
box -16 -6 32 210
use FILL  FILL_622
timestamp 1018054153
transform 1 0 4512 0 -1 7280
box -16 -6 32 210
use FILL  FILL_624
timestamp 1018054153
transform 1 0 4528 0 -1 7280
box -16 -6 32 210
use FILL  FILL_626
timestamp 1018054153
transform 1 0 4544 0 -1 7280
box -16 -6 32 210
use FILL  FILL_628
timestamp 1018054153
transform 1 0 4560 0 -1 7280
box -16 -6 32 210
use FILL  FILL_630
timestamp 1018054153
transform 1 0 4576 0 -1 7280
box -16 -6 32 210
use FILL  FILL_632
timestamp 1018054153
transform 1 0 4592 0 -1 7280
box -16 -6 32 210
use FILL  FILL_634
timestamp 1018054153
transform 1 0 4608 0 -1 7280
box -16 -6 32 210
use FILL  FILL_636
timestamp 1018054153
transform 1 0 4624 0 -1 7280
box -16 -6 32 210
use FILL  FILL_638
timestamp 1018054153
transform 1 0 4640 0 -1 7280
box -16 -6 32 210
use FILL  FILL_640
timestamp 1018054153
transform 1 0 4656 0 -1 7280
box -16 -6 32 210
use FILL  FILL_642
timestamp 1018054153
transform 1 0 4672 0 -1 7280
box -16 -6 32 210
use FILL  FILL_644
timestamp 1018054153
transform 1 0 4688 0 -1 7280
box -16 -6 32 210
use FILL  FILL_646
timestamp 1018054153
transform 1 0 4704 0 -1 7280
box -16 -6 32 210
use FILL  FILL_648
timestamp 1018054153
transform 1 0 4720 0 -1 7280
box -16 -6 32 210
use FILL  FILL_650
timestamp 1018054153
transform 1 0 4736 0 -1 7280
box -16 -6 32 210
use FILL  FILL_652
timestamp 1018054153
transform 1 0 4752 0 -1 7280
box -16 -6 32 210
use FILL  FILL_654
timestamp 1018054153
transform 1 0 4768 0 -1 7280
box -16 -6 32 210
use FILL  FILL_656
timestamp 1018054153
transform 1 0 4784 0 -1 7280
box -16 -6 32 210
use FILL  FILL_658
timestamp 1018054153
transform 1 0 4800 0 -1 7280
box -16 -6 32 210
use FILL  FILL_660
timestamp 1018054153
transform 1 0 4816 0 -1 7280
box -16 -6 32 210
use FILL  FILL_662
timestamp 1018054153
transform 1 0 4832 0 -1 7280
box -16 -6 32 210
use FILL  FILL_664
timestamp 1018054153
transform 1 0 4848 0 -1 7280
box -16 -6 32 210
use FILL  FILL_666
timestamp 1018054153
transform 1 0 4864 0 -1 7280
box -16 -6 32 210
use FILL  FILL_668
timestamp 1018054153
transform 1 0 4880 0 -1 7280
box -16 -6 32 210
use FILL  FILL_670
timestamp 1018054153
transform 1 0 4896 0 -1 7280
box -16 -6 32 210
use FILL  FILL_672
timestamp 1018054153
transform 1 0 4912 0 -1 7280
box -16 -6 32 210
use FILL  FILL_674
timestamp 1018054153
transform 1 0 4928 0 -1 7280
box -16 -6 32 210
use FILL  FILL_676
timestamp 1018054153
transform 1 0 4944 0 -1 7280
box -16 -6 32 210
use FILL  FILL_678
timestamp 1018054153
transform 1 0 4960 0 -1 7280
box -16 -6 32 210
use FILL  FILL_680
timestamp 1018054153
transform 1 0 4976 0 -1 7280
box -16 -6 32 210
use FILL  FILL_682
timestamp 1018054153
transform 1 0 4992 0 -1 7280
box -16 -6 32 210
use FILL  FILL_684
timestamp 1018054153
transform 1 0 5008 0 -1 7280
box -16 -6 32 210
use FILL  FILL_686
timestamp 1018054153
transform 1 0 5024 0 -1 7280
box -16 -6 32 210
use FILL  FILL_688
timestamp 1018054153
transform 1 0 5040 0 -1 7280
box -16 -6 32 210
use FILL  FILL_690
timestamp 1018054153
transform 1 0 5056 0 -1 7280
box -16 -6 32 210
use FILL  FILL_692
timestamp 1018054153
transform 1 0 5072 0 -1 7280
box -16 -6 32 210
use FILL  FILL_694
timestamp 1018054153
transform 1 0 5088 0 -1 7280
box -16 -6 32 210
use FILL  FILL_696
timestamp 1018054153
transform 1 0 5104 0 -1 7280
box -16 -6 32 210
use FILL  FILL_698
timestamp 1018054153
transform 1 0 5120 0 -1 7280
box -16 -6 32 210
use FILL  FILL_700
timestamp 1018054153
transform 1 0 5136 0 -1 7280
box -16 -6 32 210
use FILL  FILL_702
timestamp 1018054153
transform 1 0 5152 0 -1 7280
box -16 -6 32 210
use FILL  FILL_704
timestamp 1018054153
transform 1 0 5168 0 -1 7280
box -16 -6 32 210
use FILL  FILL_706
timestamp 1018054153
transform 1 0 5184 0 -1 7280
box -16 -6 32 210
use FILL  FILL_708
timestamp 1018054153
transform 1 0 5200 0 -1 7280
box -16 -6 32 210
use FILL  FILL_710
timestamp 1018054153
transform 1 0 5216 0 -1 7280
box -16 -6 32 210
use FILL  FILL_712
timestamp 1018054153
transform 1 0 5232 0 -1 7280
box -16 -6 32 210
use FILL  FILL_714
timestamp 1018054153
transform 1 0 5248 0 -1 7280
box -16 -6 32 210
use FILL  FILL_716
timestamp 1018054153
transform 1 0 5264 0 -1 7280
box -16 -6 32 210
use FILL  FILL_718
timestamp 1018054153
transform 1 0 5280 0 -1 7280
box -16 -6 32 210
use FILL  FILL_720
timestamp 1018054153
transform 1 0 5296 0 -1 7280
box -16 -6 32 210
use FILL  FILL_722
timestamp 1018054153
transform 1 0 5312 0 -1 7280
box -16 -6 32 210
use FILL  FILL_724
timestamp 1018054153
transform 1 0 5328 0 -1 7280
box -16 -6 32 210
use FILL  FILL_726
timestamp 1018054153
transform 1 0 5344 0 -1 7280
box -16 -6 32 210
use FILL  FILL_728
timestamp 1018054153
transform 1 0 5360 0 -1 7280
box -16 -6 32 210
use FILL  FILL_730
timestamp 1018054153
transform 1 0 5376 0 -1 7280
box -16 -6 32 210
use FILL  FILL_732
timestamp 1018054153
transform 1 0 5392 0 -1 7280
box -16 -6 32 210
use FILL  FILL_734
timestamp 1018054153
transform 1 0 5408 0 -1 7280
box -16 -6 32 210
use FILL  FILL_736
timestamp 1018054153
transform 1 0 5424 0 -1 7280
box -16 -6 32 210
use FILL  FILL_738
timestamp 1018054153
transform 1 0 5440 0 -1 7280
box -16 -6 32 210
use FILL  FILL_740
timestamp 1018054153
transform 1 0 5456 0 -1 7280
box -16 -6 32 210
use FILL  FILL_742
timestamp 1018054153
transform 1 0 5472 0 -1 7280
box -16 -6 32 210
use FILL  FILL_744
timestamp 1018054153
transform 1 0 5488 0 -1 7280
box -16 -6 32 210
use FILL  FILL_746
timestamp 1018054153
transform 1 0 5504 0 -1 7280
box -16 -6 32 210
use FILL  FILL_748
timestamp 1018054153
transform 1 0 5520 0 -1 7280
box -16 -6 32 210
use FILL  FILL_750
timestamp 1018054153
transform 1 0 5536 0 -1 7280
box -16 -6 32 210
use FILL  FILL_752
timestamp 1018054153
transform 1 0 5552 0 -1 7280
box -16 -6 32 210
use FILL  FILL_754
timestamp 1018054153
transform 1 0 5568 0 -1 7280
box -16 -6 32 210
use FILL  FILL_756
timestamp 1018054153
transform 1 0 5584 0 -1 7280
box -16 -6 32 210
use FILL  FILL_758
timestamp 1018054153
transform 1 0 5600 0 -1 7280
box -16 -6 32 210
use FILL  FILL_760
timestamp 1018054153
transform 1 0 5616 0 -1 7280
box -16 -6 32 210
use FILL  FILL_762
timestamp 1018054153
transform 1 0 5632 0 -1 7280
box -16 -6 32 210
use FILL  FILL_764
timestamp 1018054153
transform 1 0 5648 0 -1 7280
box -16 -6 32 210
use FILL  FILL_766
timestamp 1018054153
transform 1 0 5664 0 -1 7280
box -16 -6 32 210
use FILL  FILL_768
timestamp 1018054153
transform 1 0 5680 0 -1 7280
box -16 -6 32 210
use FILL  FILL_770
timestamp 1018054153
transform 1 0 5696 0 -1 7280
box -16 -6 32 210
use FILL  FILL_772
timestamp 1018054153
transform 1 0 5712 0 -1 7280
box -16 -6 32 210
use FILL  FILL_774
timestamp 1018054153
transform 1 0 5728 0 -1 7280
box -16 -6 32 210
use FILL  FILL_776
timestamp 1018054153
transform 1 0 5744 0 -1 7280
box -16 -6 32 210
use FILL  FILL_778
timestamp 1018054153
transform 1 0 5760 0 -1 7280
box -16 -6 32 210
use FILL  FILL_780
timestamp 1018054153
transform 1 0 5776 0 -1 7280
box -16 -6 32 210
use FILL  FILL_782
timestamp 1018054153
transform 1 0 5792 0 -1 7280
box -16 -6 32 210
use FILL  FILL_784
timestamp 1018054153
transform 1 0 5808 0 -1 7280
box -16 -6 32 210
use FILL  FILL_786
timestamp 1018054153
transform 1 0 5824 0 -1 7280
box -16 -6 32 210
use FILL  FILL_788
timestamp 1018054153
transform 1 0 5840 0 -1 7280
box -16 -6 32 210
use FILL  FILL_790
timestamp 1018054153
transform 1 0 5856 0 -1 7280
box -16 -6 32 210
use FILL  FILL_792
timestamp 1018054153
transform 1 0 5872 0 -1 7280
box -16 -6 32 210
use FILL  FILL_794
timestamp 1018054153
transform 1 0 5888 0 -1 7280
box -16 -6 32 210
use FILL  FILL_796
timestamp 1018054153
transform 1 0 5904 0 -1 7280
box -16 -6 32 210
use FILL  FILL_798
timestamp 1018054153
transform 1 0 5920 0 -1 7280
box -16 -6 32 210
use FILL  FILL_800
timestamp 1018054153
transform 1 0 5936 0 -1 7280
box -16 -6 32 210
use FILL  FILL_802
timestamp 1018054153
transform 1 0 5952 0 -1 7280
box -16 -6 32 210
use FILL  FILL_804
timestamp 1018054153
transform 1 0 5968 0 -1 7280
box -16 -6 32 210
use FILL  FILL_806
timestamp 1018054153
transform 1 0 5984 0 -1 7280
box -16 -6 32 210
use FILL  FILL_808
timestamp 1018054153
transform 1 0 6000 0 -1 7280
box -16 -6 32 210
use FILL  FILL_810
timestamp 1018054153
transform 1 0 6016 0 -1 7280
box -16 -6 32 210
use FILL  FILL_812
timestamp 1018054153
transform 1 0 6032 0 -1 7280
box -16 -6 32 210
use FILL  FILL_814
timestamp 1018054153
transform 1 0 6048 0 -1 7280
box -16 -6 32 210
use FILL  FILL_816
timestamp 1018054153
transform 1 0 6064 0 -1 7280
box -16 -6 32 210
use FILL  FILL_818
timestamp 1018054153
transform 1 0 6080 0 -1 7280
box -16 -6 32 210
use FILL  FILL_820
timestamp 1018054153
transform 1 0 6096 0 -1 7280
box -16 -6 32 210
use FILL  FILL_822
timestamp 1018054153
transform 1 0 6112 0 -1 7280
box -16 -6 32 210
use FILL  FILL_824
timestamp 1018054153
transform 1 0 6128 0 -1 7280
box -16 -6 32 210
use FILL  FILL_826
timestamp 1018054153
transform 1 0 6144 0 -1 7280
box -16 -6 32 210
use FILL  FILL_828
timestamp 1018054153
transform 1 0 6160 0 -1 7280
box -16 -6 32 210
use FILL  FILL_830
timestamp 1018054153
transform 1 0 6176 0 -1 7280
box -16 -6 32 210
use FILL  FILL_832
timestamp 1018054153
transform 1 0 6192 0 -1 7280
box -16 -6 32 210
use FILL  FILL_834
timestamp 1018054153
transform 1 0 6208 0 -1 7280
box -16 -6 32 210
use FILL  FILL_836
timestamp 1018054153
transform 1 0 6224 0 -1 7280
box -16 -6 32 210
use FILL  FILL_838
timestamp 1018054153
transform 1 0 6240 0 -1 7280
box -16 -6 32 210
use FILL  FILL_840
timestamp 1018054153
transform 1 0 6256 0 -1 7280
box -16 -6 32 210
use FILL  FILL_842
timestamp 1018054153
transform 1 0 6272 0 -1 7280
box -16 -6 32 210
use FILL  FILL_844
timestamp 1018054153
transform 1 0 6288 0 -1 7280
box -16 -6 32 210
use FILL  FILL_846
timestamp 1018054153
transform 1 0 6304 0 -1 7280
box -16 -6 32 210
use FILL  FILL_848
timestamp 1018054153
transform 1 0 6320 0 -1 7280
box -16 -6 32 210
use FILL  FILL_850
timestamp 1018054153
transform 1 0 6336 0 -1 7280
box -16 -6 32 210
use FILL  FILL_852
timestamp 1018054153
transform 1 0 6352 0 -1 7280
box -16 -6 32 210
use FILL  FILL_854
timestamp 1018054153
transform 1 0 6368 0 -1 7280
box -16 -6 32 210
use FILL  FILL_856
timestamp 1018054153
transform 1 0 6384 0 -1 7280
box -16 -6 32 210
use FILL  FILL_858
timestamp 1018054153
transform 1 0 6400 0 -1 7280
box -16 -6 32 210
use FILL  FILL_860
timestamp 1018054153
transform 1 0 6416 0 -1 7280
box -16 -6 32 210
use FILL  FILL_862
timestamp 1018054153
transform 1 0 6432 0 -1 7280
box -16 -6 32 210
use FILL  FILL_864
timestamp 1018054153
transform 1 0 6448 0 -1 7280
box -16 -6 32 210
use FILL  FILL_866
timestamp 1018054153
transform 1 0 6464 0 -1 7280
box -16 -6 32 210
use FILL  FILL_868
timestamp 1018054153
transform 1 0 6480 0 -1 7280
box -16 -6 32 210
use FILL  FILL_870
timestamp 1018054153
transform 1 0 6496 0 -1 7280
box -16 -6 32 210
use FILL  FILL_872
timestamp 1018054153
transform 1 0 6512 0 -1 7280
box -16 -6 32 210
use FILL  FILL_874
timestamp 1018054153
transform 1 0 6528 0 -1 7280
box -16 -6 32 210
use FILL  FILL_876
timestamp 1018054153
transform 1 0 6544 0 -1 7280
box -16 -6 32 210
use FILL  FILL_878
timestamp 1018054153
transform 1 0 6560 0 -1 7280
box -16 -6 32 210
use FILL  FILL_880
timestamp 1018054153
transform 1 0 6576 0 -1 7280
box -16 -6 32 210
use FILL  FILL_882
timestamp 1018054153
transform 1 0 6592 0 -1 7280
box -16 -6 32 210
use FILL  FILL_884
timestamp 1018054153
transform 1 0 6608 0 -1 7280
box -16 -6 32 210
use FILL  FILL_886
timestamp 1018054153
transform 1 0 6624 0 -1 7280
box -16 -6 32 210
use FILL  FILL_888
timestamp 1018054153
transform 1 0 6640 0 -1 7280
box -16 -6 32 210
use FILL  FILL_890
timestamp 1018054153
transform 1 0 6656 0 -1 7280
box -16 -6 32 210
use FILL  FILL_892
timestamp 1018054153
transform 1 0 6672 0 -1 7280
box -16 -6 32 210
use FILL  FILL_894
timestamp 1018054153
transform 1 0 6688 0 -1 7280
box -16 -6 32 210
use FILL  FILL_896
timestamp 1018054153
transform 1 0 6704 0 -1 7280
box -16 -6 32 210
use FILL  FILL_898
timestamp 1018054153
transform 1 0 6720 0 -1 7280
box -16 -6 32 210
use FILL  FILL_900
timestamp 1018054153
transform 1 0 6736 0 -1 7280
box -16 -6 32 210
use FILL  FILL_902
timestamp 1018054153
transform 1 0 6752 0 -1 7280
box -16 -6 32 210
use FILL  FILL_904
timestamp 1018054153
transform 1 0 6768 0 -1 7280
box -16 -6 32 210
use FILL  FILL_906
timestamp 1018054153
transform 1 0 6784 0 -1 7280
box -16 -6 32 210
use FILL  FILL_908
timestamp 1018054153
transform 1 0 6800 0 -1 7280
box -16 -6 32 210
use FILL  FILL_910
timestamp 1018054153
transform 1 0 6816 0 -1 7280
box -16 -6 32 210
use FILL  FILL_912
timestamp 1018054153
transform 1 0 6832 0 -1 7280
box -16 -6 32 210
use FILL  FILL_914
timestamp 1018054153
transform 1 0 6848 0 -1 7280
box -16 -6 32 210
use FILL  FILL_916
timestamp 1018054153
transform 1 0 6864 0 -1 7280
box -16 -6 32 210
use FILL  FILL_918
timestamp 1018054153
transform 1 0 6880 0 -1 7280
box -16 -6 32 210
use FILL  FILL_920
timestamp 1018054153
transform 1 0 6896 0 -1 7280
box -16 -6 32 210
use FILL  FILL_922
timestamp 1018054153
transform 1 0 6912 0 -1 7280
box -16 -6 32 210
use FILL  FILL_924
timestamp 1018054153
transform 1 0 6928 0 -1 7280
box -16 -6 32 210
use FILL  FILL_926
timestamp 1018054153
transform 1 0 6944 0 -1 7280
box -16 -6 32 210
use FILL  FILL_928
timestamp 1018054153
transform 1 0 6960 0 -1 7280
box -16 -6 32 210
use FILL  FILL_930
timestamp 1018054153
transform 1 0 6976 0 -1 7280
box -16 -6 32 210
use FILL  FILL_932
timestamp 1018054153
transform 1 0 6992 0 -1 7280
box -16 -6 32 210
use FILL  FILL_934
timestamp 1018054153
transform 1 0 7008 0 -1 7280
box -16 -6 32 210
use FILL  FILL_936
timestamp 1018054153
transform 1 0 7024 0 -1 7280
box -16 -6 32 210
use FILL  FILL_938
timestamp 1018054153
transform 1 0 7040 0 -1 7280
box -16 -6 32 210
use FILL  FILL_940
timestamp 1018054153
transform 1 0 7056 0 -1 7280
box -16 -6 32 210
use FILL  FILL_942
timestamp 1018054153
transform 1 0 7072 0 -1 7280
box -16 -6 32 210
use FILL  FILL_944
timestamp 1018054153
transform 1 0 7088 0 -1 7280
box -16 -6 32 210
use FILL  FILL_946
timestamp 1018054153
transform 1 0 7104 0 -1 7280
box -16 -6 32 210
use FILL  FILL_948
timestamp 1018054153
transform 1 0 7120 0 -1 7280
box -16 -6 32 210
use FILL  FILL_950
timestamp 1018054153
transform 1 0 7136 0 -1 7280
box -16 -6 32 210
use FILL  FILL_952
timestamp 1018054153
transform 1 0 7152 0 -1 7280
box -16 -6 32 210
use FILL  FILL_954
timestamp 1018054153
transform 1 0 7168 0 -1 7280
box -16 -6 32 210
use FILL  FILL_956
timestamp 1018054153
transform 1 0 7184 0 -1 7280
box -16 -6 32 210
use FILL  FILL_958
timestamp 1018054153
transform 1 0 7200 0 -1 7280
box -16 -6 32 210
use FILL  FILL_960
timestamp 1018054153
transform 1 0 7216 0 -1 7280
box -16 -6 32 210
use FILL  FILL_962
timestamp 1018054153
transform 1 0 7232 0 -1 7280
box -16 -6 32 210
use FILL  FILL_964
timestamp 1018054153
transform 1 0 7248 0 -1 7280
box -16 -6 32 210
use FILL  FILL_966
timestamp 1018054153
transform 1 0 7264 0 -1 7280
box -16 -6 32 210
use FILL  FILL_968
timestamp 1018054153
transform 1 0 7280 0 -1 7280
box -16 -6 32 210
use FILL  FILL_970
timestamp 1018054153
transform 1 0 7296 0 -1 7280
box -16 -6 32 210
use FILL  FILL_972
timestamp 1018054153
transform 1 0 7312 0 -1 7280
box -16 -6 32 210
use FILL  FILL_974
timestamp 1018054153
transform 1 0 7328 0 -1 7280
box -16 -6 32 210
use FILL  FILL_976
timestamp 1018054153
transform 1 0 7344 0 -1 7280
box -16 -6 32 210
use FILL  FILL_978
timestamp 1018054153
transform 1 0 7360 0 -1 7280
box -16 -6 32 210
use FILL  FILL_980
timestamp 1018054153
transform 1 0 7376 0 -1 7280
box -16 -6 32 210
use FILL  FILL_982
timestamp 1018054153
transform 1 0 7392 0 -1 7280
box -16 -6 32 210
use FILL  FILL_984
timestamp 1018054153
transform 1 0 7408 0 -1 7280
box -16 -6 32 210
use FILL  FILL_986
timestamp 1018054153
transform 1 0 7424 0 -1 7280
box -16 -6 32 210
use FILL  FILL_988
timestamp 1018054153
transform 1 0 7440 0 -1 7280
box -16 -6 32 210
use FILL  FILL_990
timestamp 1018054153
transform 1 0 7456 0 -1 7280
box -16 -6 32 210
use FILL  FILL_992
timestamp 1018054153
transform 1 0 7472 0 -1 7280
box -16 -6 32 210
use FILL  FILL_994
timestamp 1018054153
transform 1 0 7488 0 -1 7280
box -16 -6 32 210
use FILL  FILL_996
timestamp 1018054153
transform 1 0 7504 0 -1 7280
box -16 -6 32 210
use FILL  FILL_998
timestamp 1018054153
transform 1 0 7520 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1000
timestamp 1018054153
transform 1 0 7536 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1002
timestamp 1018054153
transform 1 0 7552 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1004
timestamp 1018054153
transform 1 0 7568 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1006
timestamp 1018054153
transform 1 0 7584 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1008
timestamp 1018054153
transform 1 0 7600 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1010
timestamp 1018054153
transform 1 0 7616 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1012
timestamp 1018054153
transform 1 0 7632 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1014
timestamp 1018054153
transform 1 0 7648 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1016
timestamp 1018054153
transform 1 0 7664 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1018
timestamp 1018054153
transform 1 0 7680 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1020
timestamp 1018054153
transform 1 0 7696 0 -1 7280
box -16 -6 32 210
use FILL  FILL_1022
timestamp 1018054153
transform 1 0 7712 0 -1 7280
box -16 -6 32 210
use mult_pad_VIA6  mult_pad_VIA6_2
timestamp 1542725905
transform 1 0 2212 0 1 7100
box -48 -96 48 96
use M2_M1  M2_M1_5
timestamp 1542725905
transform 1 0 4328 0 1 6950
box -4 -4 4 4
use M2_M1  M2_M1_3
timestamp 1542725905
transform 1 0 4408 0 1 6990
box -4 -4 4 4
use M2_M1  M2_M1_4
timestamp 1542725905
transform 1 0 4408 0 1 6970
box -4 -4 4 4
use M2_M1  M2_M1_2
timestamp 1542725905
transform 1 0 4552 0 1 7010
box -4 -4 4 4
use M2_M1  M2_M1_6
timestamp 1542725905
transform 1 0 5128 0 1 6950
box -4 -4 4 4
use M2_M1  M2_M1_7
timestamp 1542725905
transform 1 0 5224 0 1 6930
box -4 -4 4 4
use M3_M2  M3_M2_1
timestamp 1542725905
transform 1 0 5240 0 1 6930
box -6 -6 6 6
use M3_M2  M3_M2_0
timestamp 1542725905
transform 1 0 6120 0 1 6950
box -6 -6 6 6
use mult_pad_VIA6  mult_pad_VIA6_3
timestamp 1542725905
transform 1 0 7788 0 1 7100
box -48 -96 48 96
use mult_pad_VIA1  mult_pad_VIA1_4
timestamp 1542725905
transform 1 0 2092 0 1 6880
box -48 -6 48 6
use FILL  FILL_1023
timestamp 1018054153
transform 1 0 2272 0 1 6880
box -16 -6 32 210
use FILL  FILL_1025
timestamp 1018054153
transform 1 0 2288 0 1 6880
box -16 -6 32 210
use FILL  FILL_1027
timestamp 1018054153
transform 1 0 2304 0 1 6880
box -16 -6 32 210
use FILL  FILL_1029
timestamp 1018054153
transform 1 0 2320 0 1 6880
box -16 -6 32 210
use FILL  FILL_1031
timestamp 1018054153
transform 1 0 2336 0 1 6880
box -16 -6 32 210
use FILL  FILL_1033
timestamp 1018054153
transform 1 0 2352 0 1 6880
box -16 -6 32 210
use FILL  FILL_1035
timestamp 1018054153
transform 1 0 2368 0 1 6880
box -16 -6 32 210
use FILL  FILL_1037
timestamp 1018054153
transform 1 0 2384 0 1 6880
box -16 -6 32 210
use FILL  FILL_1039
timestamp 1018054153
transform 1 0 2400 0 1 6880
box -16 -6 32 210
use FILL  FILL_1041
timestamp 1018054153
transform 1 0 2416 0 1 6880
box -16 -6 32 210
use FILL  FILL_1043
timestamp 1018054153
transform 1 0 2432 0 1 6880
box -16 -6 32 210
use FILL  FILL_1045
timestamp 1018054153
transform 1 0 2448 0 1 6880
box -16 -6 32 210
use FILL  FILL_1047
timestamp 1018054153
transform 1 0 2464 0 1 6880
box -16 -6 32 210
use FILL  FILL_1049
timestamp 1018054153
transform 1 0 2480 0 1 6880
box -16 -6 32 210
use FILL  FILL_1051
timestamp 1018054153
transform 1 0 2496 0 1 6880
box -16 -6 32 210
use FILL  FILL_1053
timestamp 1018054153
transform 1 0 2512 0 1 6880
box -16 -6 32 210
use FILL  FILL_1055
timestamp 1018054153
transform 1 0 2528 0 1 6880
box -16 -6 32 210
use FILL  FILL_1057
timestamp 1018054153
transform 1 0 2544 0 1 6880
box -16 -6 32 210
use FILL  FILL_1059
timestamp 1018054153
transform 1 0 2560 0 1 6880
box -16 -6 32 210
use FILL  FILL_1061
timestamp 1018054153
transform 1 0 2576 0 1 6880
box -16 -6 32 210
use FILL  FILL_1063
timestamp 1018054153
transform 1 0 2592 0 1 6880
box -16 -6 32 210
use FILL  FILL_1065
timestamp 1018054153
transform 1 0 2608 0 1 6880
box -16 -6 32 210
use FILL  FILL_1067
timestamp 1018054153
transform 1 0 2624 0 1 6880
box -16 -6 32 210
use FILL  FILL_1069
timestamp 1018054153
transform 1 0 2640 0 1 6880
box -16 -6 32 210
use FILL  FILL_1071
timestamp 1018054153
transform 1 0 2656 0 1 6880
box -16 -6 32 210
use FILL  FILL_1073
timestamp 1018054153
transform 1 0 2672 0 1 6880
box -16 -6 32 210
use FILL  FILL_1075
timestamp 1018054153
transform 1 0 2688 0 1 6880
box -16 -6 32 210
use FILL  FILL_1077
timestamp 1018054153
transform 1 0 2704 0 1 6880
box -16 -6 32 210
use FILL  FILL_1079
timestamp 1018054153
transform 1 0 2720 0 1 6880
box -16 -6 32 210
use FILL  FILL_1081
timestamp 1018054153
transform 1 0 2736 0 1 6880
box -16 -6 32 210
use FILL  FILL_1083
timestamp 1018054153
transform 1 0 2752 0 1 6880
box -16 -6 32 210
use FILL  FILL_1085
timestamp 1018054153
transform 1 0 2768 0 1 6880
box -16 -6 32 210
use FILL  FILL_1087
timestamp 1018054153
transform 1 0 2784 0 1 6880
box -16 -6 32 210
use FILL  FILL_1089
timestamp 1018054153
transform 1 0 2800 0 1 6880
box -16 -6 32 210
use FILL  FILL_1091
timestamp 1018054153
transform 1 0 2816 0 1 6880
box -16 -6 32 210
use FILL  FILL_1093
timestamp 1018054153
transform 1 0 2832 0 1 6880
box -16 -6 32 210
use FILL  FILL_1095
timestamp 1018054153
transform 1 0 2848 0 1 6880
box -16 -6 32 210
use FILL  FILL_1097
timestamp 1018054153
transform 1 0 2864 0 1 6880
box -16 -6 32 210
use FILL  FILL_1099
timestamp 1018054153
transform 1 0 2880 0 1 6880
box -16 -6 32 210
use FILL  FILL_1101
timestamp 1018054153
transform 1 0 2896 0 1 6880
box -16 -6 32 210
use FILL  FILL_1103
timestamp 1018054153
transform 1 0 2912 0 1 6880
box -16 -6 32 210
use FILL  FILL_1105
timestamp 1018054153
transform 1 0 2928 0 1 6880
box -16 -6 32 210
use FILL  FILL_1107
timestamp 1018054153
transform 1 0 2944 0 1 6880
box -16 -6 32 210
use FILL  FILL_1109
timestamp 1018054153
transform 1 0 2960 0 1 6880
box -16 -6 32 210
use FILL  FILL_1111
timestamp 1018054153
transform 1 0 2976 0 1 6880
box -16 -6 32 210
use FILL  FILL_1113
timestamp 1018054153
transform 1 0 2992 0 1 6880
box -16 -6 32 210
use FILL  FILL_1115
timestamp 1018054153
transform 1 0 3008 0 1 6880
box -16 -6 32 210
use FILL  FILL_1117
timestamp 1018054153
transform 1 0 3024 0 1 6880
box -16 -6 32 210
use FILL  FILL_1119
timestamp 1018054153
transform 1 0 3040 0 1 6880
box -16 -6 32 210
use FILL  FILL_1121
timestamp 1018054153
transform 1 0 3056 0 1 6880
box -16 -6 32 210
use FILL  FILL_1123
timestamp 1018054153
transform 1 0 3072 0 1 6880
box -16 -6 32 210
use FILL  FILL_1125
timestamp 1018054153
transform 1 0 3088 0 1 6880
box -16 -6 32 210
use FILL  FILL_1127
timestamp 1018054153
transform 1 0 3104 0 1 6880
box -16 -6 32 210
use FILL  FILL_1129
timestamp 1018054153
transform 1 0 3120 0 1 6880
box -16 -6 32 210
use FILL  FILL_1131
timestamp 1018054153
transform 1 0 3136 0 1 6880
box -16 -6 32 210
use FILL  FILL_1133
timestamp 1018054153
transform 1 0 3152 0 1 6880
box -16 -6 32 210
use FILL  FILL_1135
timestamp 1018054153
transform 1 0 3168 0 1 6880
box -16 -6 32 210
use FILL  FILL_1137
timestamp 1018054153
transform 1 0 3184 0 1 6880
box -16 -6 32 210
use FILL  FILL_1139
timestamp 1018054153
transform 1 0 3200 0 1 6880
box -16 -6 32 210
use FILL  FILL_1141
timestamp 1018054153
transform 1 0 3216 0 1 6880
box -16 -6 32 210
use FILL  FILL_1143
timestamp 1018054153
transform 1 0 3232 0 1 6880
box -16 -6 32 210
use FILL  FILL_1145
timestamp 1018054153
transform 1 0 3248 0 1 6880
box -16 -6 32 210
use FILL  FILL_1147
timestamp 1018054153
transform 1 0 3264 0 1 6880
box -16 -6 32 210
use FILL  FILL_1149
timestamp 1018054153
transform 1 0 3280 0 1 6880
box -16 -6 32 210
use FILL  FILL_1151
timestamp 1018054153
transform 1 0 3296 0 1 6880
box -16 -6 32 210
use FILL  FILL_1153
timestamp 1018054153
transform 1 0 3312 0 1 6880
box -16 -6 32 210
use FILL  FILL_1155
timestamp 1018054153
transform 1 0 3328 0 1 6880
box -16 -6 32 210
use FILL  FILL_1157
timestamp 1018054153
transform 1 0 3344 0 1 6880
box -16 -6 32 210
use FILL  FILL_1159
timestamp 1018054153
transform 1 0 3360 0 1 6880
box -16 -6 32 210
use FILL  FILL_1161
timestamp 1018054153
transform 1 0 3376 0 1 6880
box -16 -6 32 210
use FILL  FILL_1163
timestamp 1018054153
transform 1 0 3392 0 1 6880
box -16 -6 32 210
use FILL  FILL_1165
timestamp 1018054153
transform 1 0 3408 0 1 6880
box -16 -6 32 210
use FILL  FILL_1167
timestamp 1018054153
transform 1 0 3424 0 1 6880
box -16 -6 32 210
use FILL  FILL_1169
timestamp 1018054153
transform 1 0 3440 0 1 6880
box -16 -6 32 210
use FILL  FILL_1171
timestamp 1018054153
transform 1 0 3456 0 1 6880
box -16 -6 32 210
use FILL  FILL_1173
timestamp 1018054153
transform 1 0 3472 0 1 6880
box -16 -6 32 210
use FILL  FILL_1175
timestamp 1018054153
transform 1 0 3488 0 1 6880
box -16 -6 32 210
use FILL  FILL_1177
timestamp 1018054153
transform 1 0 3504 0 1 6880
box -16 -6 32 210
use FILL  FILL_1179
timestamp 1018054153
transform 1 0 3520 0 1 6880
box -16 -6 32 210
use FILL  FILL_1181
timestamp 1018054153
transform 1 0 3536 0 1 6880
box -16 -6 32 210
use FILL  FILL_1183
timestamp 1018054153
transform 1 0 3552 0 1 6880
box -16 -6 32 210
use FILL  FILL_1185
timestamp 1018054153
transform 1 0 3568 0 1 6880
box -16 -6 32 210
use FILL  FILL_1187
timestamp 1018054153
transform 1 0 3584 0 1 6880
box -16 -6 32 210
use FILL  FILL_1189
timestamp 1018054153
transform 1 0 3600 0 1 6880
box -16 -6 32 210
use FILL  FILL_1191
timestamp 1018054153
transform 1 0 3616 0 1 6880
box -16 -6 32 210
use FILL  FILL_1193
timestamp 1018054153
transform 1 0 3632 0 1 6880
box -16 -6 32 210
use FILL  FILL_1195
timestamp 1018054153
transform 1 0 3648 0 1 6880
box -16 -6 32 210
use FILL  FILL_1197
timestamp 1018054153
transform 1 0 3664 0 1 6880
box -16 -6 32 210
use FILL  FILL_1199
timestamp 1018054153
transform 1 0 3680 0 1 6880
box -16 -6 32 210
use FILL  FILL_1201
timestamp 1018054153
transform 1 0 3696 0 1 6880
box -16 -6 32 210
use FILL  FILL_1203
timestamp 1018054153
transform 1 0 3712 0 1 6880
box -16 -6 32 210
use FILL  FILL_1205
timestamp 1018054153
transform 1 0 3728 0 1 6880
box -16 -6 32 210
use FILL  FILL_1207
timestamp 1018054153
transform 1 0 3744 0 1 6880
box -16 -6 32 210
use FILL  FILL_1209
timestamp 1018054153
transform 1 0 3760 0 1 6880
box -16 -6 32 210
use FILL  FILL_1211
timestamp 1018054153
transform 1 0 3776 0 1 6880
box -16 -6 32 210
use FILL  FILL_1213
timestamp 1018054153
transform 1 0 3792 0 1 6880
box -16 -6 32 210
use FILL  FILL_1215
timestamp 1018054153
transform 1 0 3808 0 1 6880
box -16 -6 32 210
use FILL  FILL_1217
timestamp 1018054153
transform 1 0 3824 0 1 6880
box -16 -6 32 210
use FILL  FILL_1219
timestamp 1018054153
transform 1 0 3840 0 1 6880
box -16 -6 32 210
use FILL  FILL_1221
timestamp 1018054153
transform 1 0 3856 0 1 6880
box -16 -6 32 210
use FILL  FILL_1223
timestamp 1018054153
transform 1 0 3872 0 1 6880
box -16 -6 32 210
use FILL  FILL_1225
timestamp 1018054153
transform 1 0 3888 0 1 6880
box -16 -6 32 210
use FILL  FILL_1227
timestamp 1018054153
transform 1 0 3904 0 1 6880
box -16 -6 32 210
use FILL  FILL_1229
timestamp 1018054153
transform 1 0 3920 0 1 6880
box -16 -6 32 210
use FILL  FILL_1231
timestamp 1018054153
transform 1 0 3936 0 1 6880
box -16 -6 32 210
use FILL  FILL_1233
timestamp 1018054153
transform 1 0 3952 0 1 6880
box -16 -6 32 210
use FILL  FILL_1235
timestamp 1018054153
transform 1 0 3968 0 1 6880
box -16 -6 32 210
use FILL  FILL_1237
timestamp 1018054153
transform 1 0 3984 0 1 6880
box -16 -6 32 210
use FILL  FILL_1239
timestamp 1018054153
transform 1 0 4000 0 1 6880
box -16 -6 32 210
use FILL  FILL_1241
timestamp 1018054153
transform 1 0 4016 0 1 6880
box -16 -6 32 210
use FILL  FILL_1243
timestamp 1018054153
transform 1 0 4032 0 1 6880
box -16 -6 32 210
use FILL  FILL_1245
timestamp 1018054153
transform 1 0 4048 0 1 6880
box -16 -6 32 210
use FILL  FILL_1247
timestamp 1018054153
transform 1 0 4064 0 1 6880
box -16 -6 32 210
use FILL  FILL_1249
timestamp 1018054153
transform 1 0 4080 0 1 6880
box -16 -6 32 210
use FILL  FILL_1251
timestamp 1018054153
transform 1 0 4096 0 1 6880
box -16 -6 32 210
use FILL  FILL_1253
timestamp 1018054153
transform 1 0 4112 0 1 6880
box -16 -6 32 210
use FILL  FILL_1255
timestamp 1018054153
transform 1 0 4128 0 1 6880
box -16 -6 32 210
use FILL  FILL_1257
timestamp 1018054153
transform 1 0 4144 0 1 6880
box -16 -6 32 210
use FILL  FILL_1259
timestamp 1018054153
transform 1 0 4160 0 1 6880
box -16 -6 32 210
use FILL  FILL_1261
timestamp 1018054153
transform 1 0 4176 0 1 6880
box -16 -6 32 210
use FILL  FILL_1263
timestamp 1018054153
transform 1 0 4192 0 1 6880
box -16 -6 32 210
use FILL  FILL_1265
timestamp 1018054153
transform 1 0 4208 0 1 6880
box -16 -6 32 210
use FILL  FILL_1267
timestamp 1018054153
transform 1 0 4224 0 1 6880
box -16 -6 32 210
use FILL  FILL_1269
timestamp 1018054153
transform 1 0 4240 0 1 6880
box -16 -6 32 210
use FILL  FILL_1271
timestamp 1018054153
transform 1 0 4256 0 1 6880
box -16 -6 32 210
use FILL  FILL_1273
timestamp 1018054153
transform 1 0 4272 0 1 6880
box -16 -6 32 210
use FILL  FILL_1275
timestamp 1018054153
transform 1 0 4288 0 1 6880
box -16 -6 32 210
use FILL  FILL_1277
timestamp 1018054153
transform 1 0 4304 0 1 6880
box -16 -6 32 210
use FILL  FILL_1279
timestamp 1018054153
transform 1 0 4320 0 1 6880
box -16 -6 32 210
use FILL  FILL_1281
timestamp 1018054153
transform 1 0 4336 0 1 6880
box -16 -6 32 210
use FILL  FILL_1282
timestamp 1018054153
transform 1 0 4352 0 1 6880
box -16 -6 32 210
use NAND2X1  NAND2X1_0
timestamp 1053022145
transform 1 0 4368 0 1 6880
box -16 -6 64 210
use FILL  FILL_1283
timestamp 1018054153
transform 1 0 4416 0 1 6880
box -16 -6 32 210
use FILL  FILL_1286
timestamp 1018054153
transform 1 0 4432 0 1 6880
box -16 -6 32 210
use FILL  FILL_1288
timestamp 1018054153
transform 1 0 4448 0 1 6880
box -16 -6 32 210
use FILL  FILL_1290
timestamp 1018054153
transform 1 0 4464 0 1 6880
box -16 -6 32 210
use FILL  FILL_1292
timestamp 1018054153
transform 1 0 4480 0 1 6880
box -16 -6 32 210
use FILL  FILL_1294
timestamp 1018054153
transform 1 0 4496 0 1 6880
box -16 -6 32 210
use FILL  FILL_1296
timestamp 1018054153
transform 1 0 4512 0 1 6880
box -16 -6 32 210
use FILL  FILL_1298
timestamp 1018054153
transform 1 0 4528 0 1 6880
box -16 -6 32 210
use FILL  FILL_1300
timestamp 1018054153
transform 1 0 4544 0 1 6880
box -16 -6 32 210
use FILL  FILL_1302
timestamp 1018054153
transform 1 0 4560 0 1 6880
box -16 -6 32 210
use FILL  FILL_1304
timestamp 1018054153
transform 1 0 4576 0 1 6880
box -16 -6 32 210
use FILL  FILL_1306
timestamp 1018054153
transform 1 0 4592 0 1 6880
box -16 -6 32 210
use FILL  FILL_1308
timestamp 1018054153
transform 1 0 4608 0 1 6880
box -16 -6 32 210
use FILL  FILL_1310
timestamp 1018054153
transform 1 0 4624 0 1 6880
box -16 -6 32 210
use FILL  FILL_1312
timestamp 1018054153
transform 1 0 4640 0 1 6880
box -16 -6 32 210
use FILL  FILL_1314
timestamp 1018054153
transform 1 0 4656 0 1 6880
box -16 -6 32 210
use FILL  FILL_1316
timestamp 1018054153
transform 1 0 4672 0 1 6880
box -16 -6 32 210
use FILL  FILL_1318
timestamp 1018054153
transform 1 0 4688 0 1 6880
box -16 -6 32 210
use FILL  FILL_1320
timestamp 1018054153
transform 1 0 4704 0 1 6880
box -16 -6 32 210
use FILL  FILL_1322
timestamp 1018054153
transform 1 0 4720 0 1 6880
box -16 -6 32 210
use FILL  FILL_1324
timestamp 1018054153
transform 1 0 4736 0 1 6880
box -16 -6 32 210
use FILL  FILL_1326
timestamp 1018054153
transform 1 0 4752 0 1 6880
box -16 -6 32 210
use FILL  FILL_1328
timestamp 1018054153
transform 1 0 4768 0 1 6880
box -16 -6 32 210
use FILL  FILL_1330
timestamp 1018054153
transform 1 0 4784 0 1 6880
box -16 -6 32 210
use FILL  FILL_1332
timestamp 1018054153
transform 1 0 4800 0 1 6880
box -16 -6 32 210
use NAND2X1  NAND2X1_1
timestamp 1053022145
transform -1 0 4864 0 1 6880
box -16 -6 64 210
use FILL  FILL_1333
timestamp 1018054153
transform 1 0 4864 0 1 6880
box -16 -6 32 210
use FILL  FILL_1337
timestamp 1018054153
transform 1 0 4880 0 1 6880
box -16 -6 32 210
use FILL  FILL_1339
timestamp 1018054153
transform 1 0 4896 0 1 6880
box -16 -6 32 210
use FILL  FILL_1341
timestamp 1018054153
transform 1 0 4912 0 1 6880
box -16 -6 32 210
use FILL  FILL_1343
timestamp 1018054153
transform 1 0 4928 0 1 6880
box -16 -6 32 210
use FILL  FILL_1345
timestamp 1018054153
transform 1 0 4944 0 1 6880
box -16 -6 32 210
use FILL  FILL_1347
timestamp 1018054153
transform 1 0 4960 0 1 6880
box -16 -6 32 210
use FILL  FILL_1349
timestamp 1018054153
transform 1 0 4976 0 1 6880
box -16 -6 32 210
use FILL  FILL_1351
timestamp 1018054153
transform 1 0 4992 0 1 6880
box -16 -6 32 210
use FILL  FILL_1353
timestamp 1018054153
transform 1 0 5008 0 1 6880
box -16 -6 32 210
use FILL  FILL_1355
timestamp 1018054153
transform 1 0 5024 0 1 6880
box -16 -6 32 210
use FILL  FILL_1357
timestamp 1018054153
transform 1 0 5040 0 1 6880
box -16 -6 32 210
use FILL  FILL_1359
timestamp 1018054153
transform 1 0 5056 0 1 6880
box -16 -6 32 210
use FILL  FILL_1361
timestamp 1018054153
transform 1 0 5072 0 1 6880
box -16 -6 32 210
use FILL  FILL_1363
timestamp 1018054153
transform 1 0 5088 0 1 6880
box -16 -6 32 210
use FILL  FILL_1365
timestamp 1018054153
transform 1 0 5104 0 1 6880
box -16 -6 32 210
use FILL  FILL_1367
timestamp 1018054153
transform 1 0 5120 0 1 6880
box -16 -6 32 210
use FILL  FILL_1369
timestamp 1018054153
transform 1 0 5136 0 1 6880
box -16 -6 32 210
use FILL  FILL_1371
timestamp 1018054153
transform 1 0 5152 0 1 6880
box -16 -6 32 210
use FILL  FILL_1373
timestamp 1018054153
transform 1 0 5168 0 1 6880
box -16 -6 32 210
use FILL  FILL_1375
timestamp 1018054153
transform 1 0 5184 0 1 6880
box -16 -6 32 210
use FILL  FILL_1376
timestamp 1018054153
transform 1 0 5200 0 1 6880
box -16 -6 32 210
use FILL  FILL_1377
timestamp 1018054153
transform 1 0 5216 0 1 6880
box -16 -6 32 210
use INVX1  INVX1_1
timestamp 1053022145
transform 1 0 5232 0 1 6880
box -18 -6 52 210
use FILL  FILL_1378
timestamp 1018054153
transform 1 0 5264 0 1 6880
box -16 -6 32 210
use FILL  FILL_1381
timestamp 1018054153
transform 1 0 5280 0 1 6880
box -16 -6 32 210
use FILL  FILL_1383
timestamp 1018054153
transform 1 0 5296 0 1 6880
box -16 -6 32 210
use FILL  FILL_1385
timestamp 1018054153
transform 1 0 5312 0 1 6880
box -16 -6 32 210
use FILL  FILL_1387
timestamp 1018054153
transform 1 0 5328 0 1 6880
box -16 -6 32 210
use FILL  FILL_1389
timestamp 1018054153
transform 1 0 5344 0 1 6880
box -16 -6 32 210
use FILL  FILL_1391
timestamp 1018054153
transform 1 0 5360 0 1 6880
box -16 -6 32 210
use FILL  FILL_1393
timestamp 1018054153
transform 1 0 5376 0 1 6880
box -16 -6 32 210
use FILL  FILL_1395
timestamp 1018054153
transform 1 0 5392 0 1 6880
box -16 -6 32 210
use FILL  FILL_1397
timestamp 1018054153
transform 1 0 5408 0 1 6880
box -16 -6 32 210
use FILL  FILL_1399
timestamp 1018054153
transform 1 0 5424 0 1 6880
box -16 -6 32 210
use FILL  FILL_1401
timestamp 1018054153
transform 1 0 5440 0 1 6880
box -16 -6 32 210
use FILL  FILL_1403
timestamp 1018054153
transform 1 0 5456 0 1 6880
box -16 -6 32 210
use FILL  FILL_1405
timestamp 1018054153
transform 1 0 5472 0 1 6880
box -16 -6 32 210
use FILL  FILL_1407
timestamp 1018054153
transform 1 0 5488 0 1 6880
box -16 -6 32 210
use FILL  FILL_1409
timestamp 1018054153
transform 1 0 5504 0 1 6880
box -16 -6 32 210
use FILL  FILL_1411
timestamp 1018054153
transform 1 0 5520 0 1 6880
box -16 -6 32 210
use FILL  FILL_1413
timestamp 1018054153
transform 1 0 5536 0 1 6880
box -16 -6 32 210
use FILL  FILL_1415
timestamp 1018054153
transform 1 0 5552 0 1 6880
box -16 -6 32 210
use FILL  FILL_1416
timestamp 1018054153
transform 1 0 5568 0 1 6880
box -16 -6 32 210
use FILL  FILL_1417
timestamp 1018054153
transform 1 0 5584 0 1 6880
box -16 -6 32 210
use FILL  FILL_1418
timestamp 1018054153
transform 1 0 5600 0 1 6880
box -16 -6 32 210
use FILL  FILL_1419
timestamp 1018054153
transform 1 0 5616 0 1 6880
box -16 -6 32 210
use FILL  FILL_1420
timestamp 1018054153
transform 1 0 5632 0 1 6880
box -16 -6 32 210
use FILL  FILL_1421
timestamp 1018054153
transform 1 0 5648 0 1 6880
box -16 -6 32 210
use FILL  FILL_1422
timestamp 1018054153
transform 1 0 5664 0 1 6880
box -16 -6 32 210
use FILL  FILL_1424
timestamp 1018054153
transform 1 0 5680 0 1 6880
box -16 -6 32 210
use FILL  FILL_1426
timestamp 1018054153
transform 1 0 5696 0 1 6880
box -16 -6 32 210
use FILL  FILL_1428
timestamp 1018054153
transform 1 0 5712 0 1 6880
box -16 -6 32 210
use FILL  FILL_1430
timestamp 1018054153
transform 1 0 5728 0 1 6880
box -16 -6 32 210
use FILL  FILL_1432
timestamp 1018054153
transform 1 0 5744 0 1 6880
box -16 -6 32 210
use FILL  FILL_1434
timestamp 1018054153
transform 1 0 5760 0 1 6880
box -16 -6 32 210
use FILL  FILL_1436
timestamp 1018054153
transform 1 0 5776 0 1 6880
box -16 -6 32 210
use FILL  FILL_1438
timestamp 1018054153
transform 1 0 5792 0 1 6880
box -16 -6 32 210
use FILL  FILL_1440
timestamp 1018054153
transform 1 0 5808 0 1 6880
box -16 -6 32 210
use FILL  FILL_1442
timestamp 1018054153
transform 1 0 5824 0 1 6880
box -16 -6 32 210
use FILL  FILL_1444
timestamp 1018054153
transform 1 0 5840 0 1 6880
box -16 -6 32 210
use FILL  FILL_1446
timestamp 1018054153
transform 1 0 5856 0 1 6880
box -16 -6 32 210
use FILL  FILL_1448
timestamp 1018054153
transform 1 0 5872 0 1 6880
box -16 -6 32 210
use FILL  FILL_1450
timestamp 1018054153
transform 1 0 5888 0 1 6880
box -16 -6 32 210
use FILL  FILL_1452
timestamp 1018054153
transform 1 0 5904 0 1 6880
box -16 -6 32 210
use FILL  FILL_1454
timestamp 1018054153
transform 1 0 5920 0 1 6880
box -16 -6 32 210
use FILL  FILL_1456
timestamp 1018054153
transform 1 0 5936 0 1 6880
box -16 -6 32 210
use FILL  FILL_1458
timestamp 1018054153
transform 1 0 5952 0 1 6880
box -16 -6 32 210
use FILL  FILL_1460
timestamp 1018054153
transform 1 0 5968 0 1 6880
box -16 -6 32 210
use FILL  FILL_1462
timestamp 1018054153
transform 1 0 5984 0 1 6880
box -16 -6 32 210
use FILL  FILL_1464
timestamp 1018054153
transform 1 0 6000 0 1 6880
box -16 -6 32 210
use FILL  FILL_1466
timestamp 1018054153
transform 1 0 6016 0 1 6880
box -16 -6 32 210
use FILL  FILL_1468
timestamp 1018054153
transform 1 0 6032 0 1 6880
box -16 -6 32 210
use FILL  FILL_1470
timestamp 1018054153
transform 1 0 6048 0 1 6880
box -16 -6 32 210
use FILL  FILL_1472
timestamp 1018054153
transform 1 0 6064 0 1 6880
box -16 -6 32 210
use FILL  FILL_1474
timestamp 1018054153
transform 1 0 6080 0 1 6880
box -16 -6 32 210
use FILL  FILL_1476
timestamp 1018054153
transform 1 0 6096 0 1 6880
box -16 -6 32 210
use FILL  FILL_1478
timestamp 1018054153
transform 1 0 6112 0 1 6880
box -16 -6 32 210
use FILL  FILL_1480
timestamp 1018054153
transform 1 0 6128 0 1 6880
box -16 -6 32 210
use FILL  FILL_1482
timestamp 1018054153
transform 1 0 6144 0 1 6880
box -16 -6 32 210
use FILL  FILL_1484
timestamp 1018054153
transform 1 0 6160 0 1 6880
box -16 -6 32 210
use FILL  FILL_1486
timestamp 1018054153
transform 1 0 6176 0 1 6880
box -16 -6 32 210
use FILL  FILL_1488
timestamp 1018054153
transform 1 0 6192 0 1 6880
box -16 -6 32 210
use FILL  FILL_1490
timestamp 1018054153
transform 1 0 6208 0 1 6880
box -16 -6 32 210
use FILL  FILL_1492
timestamp 1018054153
transform 1 0 6224 0 1 6880
box -16 -6 32 210
use FILL  FILL_1494
timestamp 1018054153
transform 1 0 6240 0 1 6880
box -16 -6 32 210
use FILL  FILL_1496
timestamp 1018054153
transform 1 0 6256 0 1 6880
box -16 -6 32 210
use FILL  FILL_1498
timestamp 1018054153
transform 1 0 6272 0 1 6880
box -16 -6 32 210
use FILL  FILL_1500
timestamp 1018054153
transform 1 0 6288 0 1 6880
box -16 -6 32 210
use FILL  FILL_1502
timestamp 1018054153
transform 1 0 6304 0 1 6880
box -16 -6 32 210
use FILL  FILL_1504
timestamp 1018054153
transform 1 0 6320 0 1 6880
box -16 -6 32 210
use FILL  FILL_1506
timestamp 1018054153
transform 1 0 6336 0 1 6880
box -16 -6 32 210
use FILL  FILL_1508
timestamp 1018054153
transform 1 0 6352 0 1 6880
box -16 -6 32 210
use FILL  FILL_1510
timestamp 1018054153
transform 1 0 6368 0 1 6880
box -16 -6 32 210
use FILL  FILL_1512
timestamp 1018054153
transform 1 0 6384 0 1 6880
box -16 -6 32 210
use FILL  FILL_1514
timestamp 1018054153
transform 1 0 6400 0 1 6880
box -16 -6 32 210
use FILL  FILL_1516
timestamp 1018054153
transform 1 0 6416 0 1 6880
box -16 -6 32 210
use FILL  FILL_1518
timestamp 1018054153
transform 1 0 6432 0 1 6880
box -16 -6 32 210
use FILL  FILL_1520
timestamp 1018054153
transform 1 0 6448 0 1 6880
box -16 -6 32 210
use FILL  FILL_1522
timestamp 1018054153
transform 1 0 6464 0 1 6880
box -16 -6 32 210
use FILL  FILL_1524
timestamp 1018054153
transform 1 0 6480 0 1 6880
box -16 -6 32 210
use FILL  FILL_1526
timestamp 1018054153
transform 1 0 6496 0 1 6880
box -16 -6 32 210
use FILL  FILL_1528
timestamp 1018054153
transform 1 0 6512 0 1 6880
box -16 -6 32 210
use FILL  FILL_1530
timestamp 1018054153
transform 1 0 6528 0 1 6880
box -16 -6 32 210
use FILL  FILL_1532
timestamp 1018054153
transform 1 0 6544 0 1 6880
box -16 -6 32 210
use FILL  FILL_1534
timestamp 1018054153
transform 1 0 6560 0 1 6880
box -16 -6 32 210
use FILL  FILL_1536
timestamp 1018054153
transform 1 0 6576 0 1 6880
box -16 -6 32 210
use FILL  FILL_1538
timestamp 1018054153
transform 1 0 6592 0 1 6880
box -16 -6 32 210
use FILL  FILL_1540
timestamp 1018054153
transform 1 0 6608 0 1 6880
box -16 -6 32 210
use FILL  FILL_1542
timestamp 1018054153
transform 1 0 6624 0 1 6880
box -16 -6 32 210
use FILL  FILL_1544
timestamp 1018054153
transform 1 0 6640 0 1 6880
box -16 -6 32 210
use FILL  FILL_1546
timestamp 1018054153
transform 1 0 6656 0 1 6880
box -16 -6 32 210
use FILL  FILL_1548
timestamp 1018054153
transform 1 0 6672 0 1 6880
box -16 -6 32 210
use FILL  FILL_1550
timestamp 1018054153
transform 1 0 6688 0 1 6880
box -16 -6 32 210
use FILL  FILL_1552
timestamp 1018054153
transform 1 0 6704 0 1 6880
box -16 -6 32 210
use FILL  FILL_1554
timestamp 1018054153
transform 1 0 6720 0 1 6880
box -16 -6 32 210
use FILL  FILL_1556
timestamp 1018054153
transform 1 0 6736 0 1 6880
box -16 -6 32 210
use FILL  FILL_1558
timestamp 1018054153
transform 1 0 6752 0 1 6880
box -16 -6 32 210
use FILL  FILL_1560
timestamp 1018054153
transform 1 0 6768 0 1 6880
box -16 -6 32 210
use FILL  FILL_1562
timestamp 1018054153
transform 1 0 6784 0 1 6880
box -16 -6 32 210
use FILL  FILL_1564
timestamp 1018054153
transform 1 0 6800 0 1 6880
box -16 -6 32 210
use FILL  FILL_1566
timestamp 1018054153
transform 1 0 6816 0 1 6880
box -16 -6 32 210
use FILL  FILL_1568
timestamp 1018054153
transform 1 0 6832 0 1 6880
box -16 -6 32 210
use FILL  FILL_1570
timestamp 1018054153
transform 1 0 6848 0 1 6880
box -16 -6 32 210
use FILL  FILL_1572
timestamp 1018054153
transform 1 0 6864 0 1 6880
box -16 -6 32 210
use FILL  FILL_1574
timestamp 1018054153
transform 1 0 6880 0 1 6880
box -16 -6 32 210
use FILL  FILL_1576
timestamp 1018054153
transform 1 0 6896 0 1 6880
box -16 -6 32 210
use FILL  FILL_1578
timestamp 1018054153
transform 1 0 6912 0 1 6880
box -16 -6 32 210
use FILL  FILL_1580
timestamp 1018054153
transform 1 0 6928 0 1 6880
box -16 -6 32 210
use FILL  FILL_1582
timestamp 1018054153
transform 1 0 6944 0 1 6880
box -16 -6 32 210
use FILL  FILL_1584
timestamp 1018054153
transform 1 0 6960 0 1 6880
box -16 -6 32 210
use FILL  FILL_1586
timestamp 1018054153
transform 1 0 6976 0 1 6880
box -16 -6 32 210
use FILL  FILL_1588
timestamp 1018054153
transform 1 0 6992 0 1 6880
box -16 -6 32 210
use FILL  FILL_1590
timestamp 1018054153
transform 1 0 7008 0 1 6880
box -16 -6 32 210
use FILL  FILL_1592
timestamp 1018054153
transform 1 0 7024 0 1 6880
box -16 -6 32 210
use FILL  FILL_1594
timestamp 1018054153
transform 1 0 7040 0 1 6880
box -16 -6 32 210
use FILL  FILL_1596
timestamp 1018054153
transform 1 0 7056 0 1 6880
box -16 -6 32 210
use FILL  FILL_1598
timestamp 1018054153
transform 1 0 7072 0 1 6880
box -16 -6 32 210
use FILL  FILL_1600
timestamp 1018054153
transform 1 0 7088 0 1 6880
box -16 -6 32 210
use FILL  FILL_1602
timestamp 1018054153
transform 1 0 7104 0 1 6880
box -16 -6 32 210
use FILL  FILL_1604
timestamp 1018054153
transform 1 0 7120 0 1 6880
box -16 -6 32 210
use FILL  FILL_1606
timestamp 1018054153
transform 1 0 7136 0 1 6880
box -16 -6 32 210
use FILL  FILL_1608
timestamp 1018054153
transform 1 0 7152 0 1 6880
box -16 -6 32 210
use FILL  FILL_1610
timestamp 1018054153
transform 1 0 7168 0 1 6880
box -16 -6 32 210
use FILL  FILL_1612
timestamp 1018054153
transform 1 0 7184 0 1 6880
box -16 -6 32 210
use FILL  FILL_1614
timestamp 1018054153
transform 1 0 7200 0 1 6880
box -16 -6 32 210
use FILL  FILL_1616
timestamp 1018054153
transform 1 0 7216 0 1 6880
box -16 -6 32 210
use FILL  FILL_1618
timestamp 1018054153
transform 1 0 7232 0 1 6880
box -16 -6 32 210
use FILL  FILL_1620
timestamp 1018054153
transform 1 0 7248 0 1 6880
box -16 -6 32 210
use FILL  FILL_1622
timestamp 1018054153
transform 1 0 7264 0 1 6880
box -16 -6 32 210
use FILL  FILL_1624
timestamp 1018054153
transform 1 0 7280 0 1 6880
box -16 -6 32 210
use FILL  FILL_1626
timestamp 1018054153
transform 1 0 7296 0 1 6880
box -16 -6 32 210
use FILL  FILL_1628
timestamp 1018054153
transform 1 0 7312 0 1 6880
box -16 -6 32 210
use FILL  FILL_1630
timestamp 1018054153
transform 1 0 7328 0 1 6880
box -16 -6 32 210
use FILL  FILL_1632
timestamp 1018054153
transform 1 0 7344 0 1 6880
box -16 -6 32 210
use FILL  FILL_1634
timestamp 1018054153
transform 1 0 7360 0 1 6880
box -16 -6 32 210
use FILL  FILL_1636
timestamp 1018054153
transform 1 0 7376 0 1 6880
box -16 -6 32 210
use FILL  FILL_1638
timestamp 1018054153
transform 1 0 7392 0 1 6880
box -16 -6 32 210
use FILL  FILL_1640
timestamp 1018054153
transform 1 0 7408 0 1 6880
box -16 -6 32 210
use FILL  FILL_1642
timestamp 1018054153
transform 1 0 7424 0 1 6880
box -16 -6 32 210
use FILL  FILL_1644
timestamp 1018054153
transform 1 0 7440 0 1 6880
box -16 -6 32 210
use FILL  FILL_1646
timestamp 1018054153
transform 1 0 7456 0 1 6880
box -16 -6 32 210
use FILL  FILL_1648
timestamp 1018054153
transform 1 0 7472 0 1 6880
box -16 -6 32 210
use FILL  FILL_1650
timestamp 1018054153
transform 1 0 7488 0 1 6880
box -16 -6 32 210
use FILL  FILL_1652
timestamp 1018054153
transform 1 0 7504 0 1 6880
box -16 -6 32 210
use FILL  FILL_1654
timestamp 1018054153
transform 1 0 7520 0 1 6880
box -16 -6 32 210
use FILL  FILL_1656
timestamp 1018054153
transform 1 0 7536 0 1 6880
box -16 -6 32 210
use FILL  FILL_1658
timestamp 1018054153
transform 1 0 7552 0 1 6880
box -16 -6 32 210
use FILL  FILL_1660
timestamp 1018054153
transform 1 0 7568 0 1 6880
box -16 -6 32 210
use FILL  FILL_1662
timestamp 1018054153
transform 1 0 7584 0 1 6880
box -16 -6 32 210
use FILL  FILL_1664
timestamp 1018054153
transform 1 0 7600 0 1 6880
box -16 -6 32 210
use FILL  FILL_1666
timestamp 1018054153
transform 1 0 7616 0 1 6880
box -16 -6 32 210
use FILL  FILL_1668
timestamp 1018054153
transform 1 0 7632 0 1 6880
box -16 -6 32 210
use FILL  FILL_1670
timestamp 1018054153
transform 1 0 7648 0 1 6880
box -16 -6 32 210
use FILL  FILL_1672
timestamp 1018054153
transform 1 0 7664 0 1 6880
box -16 -6 32 210
use FILL  FILL_1674
timestamp 1018054153
transform 1 0 7680 0 1 6880
box -16 -6 32 210
use FILL  FILL_1676
timestamp 1018054153
transform 1 0 7696 0 1 6880
box -16 -6 32 210
use FILL  FILL_1678
timestamp 1018054153
transform 1 0 7712 0 1 6880
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_5
timestamp 1542725905
transform 1 0 7908 0 1 6880
box -48 -6 48 6
use PADVDD  PADVDD_1
timestamp 1084294447
transform 0 -1 2000 1 0 6800
box -6 -6 606 2000
use M3_M2  M3_M2_2
timestamp 1542725905
transform 1 0 1998 0 1 6730
box -6 -6 6 6
use M3_M2  M3_M2_3
timestamp 1542725905
transform 1 0 4136 0 1 6730
box -6 -6 6 6
use M2_M1  M2_M1_9
timestamp 1542725905
transform 1 0 4232 0 1 6810
box -4 -4 4 4
use M2_M1  M2_M1_10
timestamp 1542725905
transform 1 0 4328 0 1 6810
box -4 -4 4 4
use M2_M1  M2_M1_11
timestamp 1542725905
transform 1 0 4392 0 1 6810
box -4 -4 4 4
use M2_M1  M2_M1_13
timestamp 1542725905
transform 1 0 4360 0 1 6790
box -4 -4 4 4
use M2_M1  M2_M1_17
timestamp 1542725905
transform 1 0 4408 0 1 6770
box -4 -4 4 4
use M2_M1  M2_M1_8
timestamp 1542725905
transform 1 0 4776 0 1 6830
box -4 -4 4 4
use M2_M1  M2_M1_12
timestamp 1542725905
transform 1 0 5160 0 1 6810
box -4 -4 4 4
use M2_M1  M2_M1_18
timestamp 1542725905
transform 1 0 5240 0 1 6770
box -4 -4 4 4
use M2_M1  M2_M1_14
timestamp 1542725905
transform 1 0 5560 0 1 6790
box -4 -4 4 4
use M2_M1  M2_M1_15
timestamp 1542725905
transform 1 0 5624 0 1 6790
box -4 -4 4 4
use M2_M1  M2_M1_16
timestamp 1542725905
transform 1 0 5704 0 1 6790
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_6
timestamp 1542725905
transform 1 0 2212 0 1 6680
box -48 -6 48 6
use FILL  FILL_1024
timestamp 1018054153
transform 1 0 2272 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1026
timestamp 1018054153
transform 1 0 2288 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1028
timestamp 1018054153
transform 1 0 2304 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1030
timestamp 1018054153
transform 1 0 2320 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1032
timestamp 1018054153
transform 1 0 2336 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1034
timestamp 1018054153
transform 1 0 2352 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1036
timestamp 1018054153
transform 1 0 2368 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1038
timestamp 1018054153
transform 1 0 2384 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1040
timestamp 1018054153
transform 1 0 2400 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1042
timestamp 1018054153
transform 1 0 2416 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1044
timestamp 1018054153
transform 1 0 2432 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1046
timestamp 1018054153
transform 1 0 2448 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1048
timestamp 1018054153
transform 1 0 2464 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1050
timestamp 1018054153
transform 1 0 2480 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1052
timestamp 1018054153
transform 1 0 2496 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1054
timestamp 1018054153
transform 1 0 2512 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1056
timestamp 1018054153
transform 1 0 2528 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1058
timestamp 1018054153
transform 1 0 2544 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1060
timestamp 1018054153
transform 1 0 2560 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1062
timestamp 1018054153
transform 1 0 2576 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1064
timestamp 1018054153
transform 1 0 2592 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1066
timestamp 1018054153
transform 1 0 2608 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1068
timestamp 1018054153
transform 1 0 2624 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1070
timestamp 1018054153
transform 1 0 2640 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1072
timestamp 1018054153
transform 1 0 2656 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1074
timestamp 1018054153
transform 1 0 2672 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1076
timestamp 1018054153
transform 1 0 2688 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1078
timestamp 1018054153
transform 1 0 2704 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1080
timestamp 1018054153
transform 1 0 2720 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1082
timestamp 1018054153
transform 1 0 2736 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1084
timestamp 1018054153
transform 1 0 2752 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1086
timestamp 1018054153
transform 1 0 2768 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1088
timestamp 1018054153
transform 1 0 2784 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1090
timestamp 1018054153
transform 1 0 2800 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1092
timestamp 1018054153
transform 1 0 2816 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1094
timestamp 1018054153
transform 1 0 2832 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1096
timestamp 1018054153
transform 1 0 2848 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1098
timestamp 1018054153
transform 1 0 2864 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1100
timestamp 1018054153
transform 1 0 2880 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1102
timestamp 1018054153
transform 1 0 2896 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1104
timestamp 1018054153
transform 1 0 2912 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1106
timestamp 1018054153
transform 1 0 2928 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1108
timestamp 1018054153
transform 1 0 2944 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1110
timestamp 1018054153
transform 1 0 2960 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1112
timestamp 1018054153
transform 1 0 2976 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1114
timestamp 1018054153
transform 1 0 2992 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1116
timestamp 1018054153
transform 1 0 3008 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1118
timestamp 1018054153
transform 1 0 3024 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1120
timestamp 1018054153
transform 1 0 3040 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1122
timestamp 1018054153
transform 1 0 3056 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1124
timestamp 1018054153
transform 1 0 3072 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1126
timestamp 1018054153
transform 1 0 3088 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1128
timestamp 1018054153
transform 1 0 3104 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1130
timestamp 1018054153
transform 1 0 3120 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1132
timestamp 1018054153
transform 1 0 3136 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1134
timestamp 1018054153
transform 1 0 3152 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1136
timestamp 1018054153
transform 1 0 3168 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1138
timestamp 1018054153
transform 1 0 3184 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1140
timestamp 1018054153
transform 1 0 3200 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1142
timestamp 1018054153
transform 1 0 3216 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1144
timestamp 1018054153
transform 1 0 3232 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1146
timestamp 1018054153
transform 1 0 3248 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1148
timestamp 1018054153
transform 1 0 3264 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1150
timestamp 1018054153
transform 1 0 3280 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1152
timestamp 1018054153
transform 1 0 3296 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1154
timestamp 1018054153
transform 1 0 3312 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1156
timestamp 1018054153
transform 1 0 3328 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1158
timestamp 1018054153
transform 1 0 3344 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1160
timestamp 1018054153
transform 1 0 3360 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1162
timestamp 1018054153
transform 1 0 3376 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1164
timestamp 1018054153
transform 1 0 3392 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1166
timestamp 1018054153
transform 1 0 3408 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1168
timestamp 1018054153
transform 1 0 3424 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1170
timestamp 1018054153
transform 1 0 3440 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1172
timestamp 1018054153
transform 1 0 3456 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1174
timestamp 1018054153
transform 1 0 3472 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1176
timestamp 1018054153
transform 1 0 3488 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1178
timestamp 1018054153
transform 1 0 3504 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1180
timestamp 1018054153
transform 1 0 3520 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1182
timestamp 1018054153
transform 1 0 3536 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1184
timestamp 1018054153
transform 1 0 3552 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1186
timestamp 1018054153
transform 1 0 3568 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1188
timestamp 1018054153
transform 1 0 3584 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1190
timestamp 1018054153
transform 1 0 3600 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1192
timestamp 1018054153
transform 1 0 3616 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1194
timestamp 1018054153
transform 1 0 3632 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1196
timestamp 1018054153
transform 1 0 3648 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1198
timestamp 1018054153
transform 1 0 3664 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1200
timestamp 1018054153
transform 1 0 3680 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1202
timestamp 1018054153
transform 1 0 3696 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1204
timestamp 1018054153
transform 1 0 3712 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1206
timestamp 1018054153
transform 1 0 3728 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1208
timestamp 1018054153
transform 1 0 3744 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1210
timestamp 1018054153
transform 1 0 3760 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1212
timestamp 1018054153
transform 1 0 3776 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1214
timestamp 1018054153
transform 1 0 3792 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1216
timestamp 1018054153
transform 1 0 3808 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1218
timestamp 1018054153
transform 1 0 3824 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1220
timestamp 1018054153
transform 1 0 3840 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1222
timestamp 1018054153
transform 1 0 3856 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1224
timestamp 1018054153
transform 1 0 3872 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1226
timestamp 1018054153
transform 1 0 3888 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1228
timestamp 1018054153
transform 1 0 3904 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1230
timestamp 1018054153
transform 1 0 3920 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1232
timestamp 1018054153
transform 1 0 3936 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1234
timestamp 1018054153
transform 1 0 3952 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1236
timestamp 1018054153
transform 1 0 3968 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1238
timestamp 1018054153
transform 1 0 3984 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1240
timestamp 1018054153
transform 1 0 4000 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1242
timestamp 1018054153
transform 1 0 4016 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1244
timestamp 1018054153
transform 1 0 4032 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1246
timestamp 1018054153
transform 1 0 4048 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1248
timestamp 1018054153
transform 1 0 4064 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1250
timestamp 1018054153
transform 1 0 4080 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1252
timestamp 1018054153
transform 1 0 4096 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1254
timestamp 1018054153
transform 1 0 4112 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1256
timestamp 1018054153
transform 1 0 4128 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1258
timestamp 1018054153
transform 1 0 4144 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1260
timestamp 1018054153
transform 1 0 4160 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1262
timestamp 1018054153
transform 1 0 4176 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1264
timestamp 1018054153
transform 1 0 4192 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1266
timestamp 1018054153
transform 1 0 4208 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1268
timestamp 1018054153
transform 1 0 4224 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1270
timestamp 1018054153
transform 1 0 4240 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1272
timestamp 1018054153
transform 1 0 4256 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1274
timestamp 1018054153
transform 1 0 4272 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1276
timestamp 1018054153
transform 1 0 4288 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1278
timestamp 1018054153
transform 1 0 4304 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1280
timestamp 1018054153
transform 1 0 4320 0 -1 6880
box -16 -6 32 210
use OAI21X1  OAI21X1_0
timestamp 1053722159
transform 1 0 4336 0 -1 6880
box -16 -6 68 210
use FILL  FILL_1284
timestamp 1018054153
transform 1 0 4400 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1285
timestamp 1018054153
transform 1 0 4416 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1287
timestamp 1018054153
transform 1 0 4432 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1289
timestamp 1018054153
transform 1 0 4448 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1291
timestamp 1018054153
transform 1 0 4464 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1293
timestamp 1018054153
transform 1 0 4480 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1295
timestamp 1018054153
transform 1 0 4496 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1297
timestamp 1018054153
transform 1 0 4512 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1299
timestamp 1018054153
transform 1 0 4528 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1301
timestamp 1018054153
transform 1 0 4544 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1303
timestamp 1018054153
transform 1 0 4560 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1305
timestamp 1018054153
transform 1 0 4576 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1307
timestamp 1018054153
transform 1 0 4592 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1309
timestamp 1018054153
transform 1 0 4608 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1311
timestamp 1018054153
transform 1 0 4624 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1313
timestamp 1018054153
transform 1 0 4640 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1315
timestamp 1018054153
transform 1 0 4656 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1317
timestamp 1018054153
transform 1 0 4672 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1319
timestamp 1018054153
transform 1 0 4688 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1321
timestamp 1018054153
transform 1 0 4704 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1323
timestamp 1018054153
transform 1 0 4720 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1325
timestamp 1018054153
transform 1 0 4736 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1327
timestamp 1018054153
transform 1 0 4752 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1329
timestamp 1018054153
transform 1 0 4768 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1331
timestamp 1018054153
transform 1 0 4784 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1334
timestamp 1018054153
transform 1 0 4800 0 -1 6880
box -16 -6 32 210
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 4816 0 -1 6880
box -18 -6 52 210
use FILL  FILL_1335
timestamp 1018054153
transform 1 0 4848 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1336
timestamp 1018054153
transform 1 0 4864 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1338
timestamp 1018054153
transform 1 0 4880 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1340
timestamp 1018054153
transform 1 0 4896 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1342
timestamp 1018054153
transform 1 0 4912 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1344
timestamp 1018054153
transform 1 0 4928 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1346
timestamp 1018054153
transform 1 0 4944 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1348
timestamp 1018054153
transform 1 0 4960 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1350
timestamp 1018054153
transform 1 0 4976 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1352
timestamp 1018054153
transform 1 0 4992 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1354
timestamp 1018054153
transform 1 0 5008 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1356
timestamp 1018054153
transform 1 0 5024 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1358
timestamp 1018054153
transform 1 0 5040 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1360
timestamp 1018054153
transform 1 0 5056 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1362
timestamp 1018054153
transform 1 0 5072 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1364
timestamp 1018054153
transform 1 0 5088 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1366
timestamp 1018054153
transform 1 0 5104 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1368
timestamp 1018054153
transform 1 0 5120 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1370
timestamp 1018054153
transform 1 0 5136 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1372
timestamp 1018054153
transform 1 0 5152 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1374
timestamp 1018054153
transform 1 0 5168 0 -1 6880
box -16 -6 32 210
use OAI21X1  OAI21X1_1
timestamp 1053722159
transform 1 0 5184 0 -1 6880
box -16 -6 68 210
use FILL  FILL_1379
timestamp 1018054153
transform 1 0 5248 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1380
timestamp 1018054153
transform 1 0 5264 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1382
timestamp 1018054153
transform 1 0 5280 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1384
timestamp 1018054153
transform 1 0 5296 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1386
timestamp 1018054153
transform 1 0 5312 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1388
timestamp 1018054153
transform 1 0 5328 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1390
timestamp 1018054153
transform 1 0 5344 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1392
timestamp 1018054153
transform 1 0 5360 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1394
timestamp 1018054153
transform 1 0 5376 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1396
timestamp 1018054153
transform 1 0 5392 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1398
timestamp 1018054153
transform 1 0 5408 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1400
timestamp 1018054153
transform 1 0 5424 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1402
timestamp 1018054153
transform 1 0 5440 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1404
timestamp 1018054153
transform 1 0 5456 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1406
timestamp 1018054153
transform 1 0 5472 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1408
timestamp 1018054153
transform 1 0 5488 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1410
timestamp 1018054153
transform 1 0 5504 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1412
timestamp 1018054153
transform 1 0 5520 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1414
timestamp 1018054153
transform 1 0 5536 0 -1 6880
box -16 -6 32 210
use XOR2X1  XOR2X1_0
timestamp 1053359338
transform 1 0 5552 0 -1 6880
box -16 -6 128 210
use FILL  FILL_1423
timestamp 1018054153
transform 1 0 5664 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1425
timestamp 1018054153
transform 1 0 5680 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1427
timestamp 1018054153
transform 1 0 5696 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1429
timestamp 1018054153
transform 1 0 5712 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1431
timestamp 1018054153
transform 1 0 5728 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1433
timestamp 1018054153
transform 1 0 5744 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1435
timestamp 1018054153
transform 1 0 5760 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1437
timestamp 1018054153
transform 1 0 5776 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1439
timestamp 1018054153
transform 1 0 5792 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1441
timestamp 1018054153
transform 1 0 5808 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1443
timestamp 1018054153
transform 1 0 5824 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1445
timestamp 1018054153
transform 1 0 5840 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1447
timestamp 1018054153
transform 1 0 5856 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1449
timestamp 1018054153
transform 1 0 5872 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1451
timestamp 1018054153
transform 1 0 5888 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1453
timestamp 1018054153
transform 1 0 5904 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1455
timestamp 1018054153
transform 1 0 5920 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1457
timestamp 1018054153
transform 1 0 5936 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1459
timestamp 1018054153
transform 1 0 5952 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1461
timestamp 1018054153
transform 1 0 5968 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1463
timestamp 1018054153
transform 1 0 5984 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1465
timestamp 1018054153
transform 1 0 6000 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1467
timestamp 1018054153
transform 1 0 6016 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1469
timestamp 1018054153
transform 1 0 6032 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1471
timestamp 1018054153
transform 1 0 6048 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1473
timestamp 1018054153
transform 1 0 6064 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1475
timestamp 1018054153
transform 1 0 6080 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1477
timestamp 1018054153
transform 1 0 6096 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1479
timestamp 1018054153
transform 1 0 6112 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1481
timestamp 1018054153
transform 1 0 6128 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1483
timestamp 1018054153
transform 1 0 6144 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1485
timestamp 1018054153
transform 1 0 6160 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1487
timestamp 1018054153
transform 1 0 6176 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1489
timestamp 1018054153
transform 1 0 6192 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1491
timestamp 1018054153
transform 1 0 6208 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1493
timestamp 1018054153
transform 1 0 6224 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1495
timestamp 1018054153
transform 1 0 6240 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1497
timestamp 1018054153
transform 1 0 6256 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1499
timestamp 1018054153
transform 1 0 6272 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1501
timestamp 1018054153
transform 1 0 6288 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1503
timestamp 1018054153
transform 1 0 6304 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1505
timestamp 1018054153
transform 1 0 6320 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1507
timestamp 1018054153
transform 1 0 6336 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1509
timestamp 1018054153
transform 1 0 6352 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1511
timestamp 1018054153
transform 1 0 6368 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1513
timestamp 1018054153
transform 1 0 6384 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1515
timestamp 1018054153
transform 1 0 6400 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1517
timestamp 1018054153
transform 1 0 6416 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1519
timestamp 1018054153
transform 1 0 6432 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1521
timestamp 1018054153
transform 1 0 6448 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1523
timestamp 1018054153
transform 1 0 6464 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1525
timestamp 1018054153
transform 1 0 6480 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1527
timestamp 1018054153
transform 1 0 6496 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1529
timestamp 1018054153
transform 1 0 6512 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1531
timestamp 1018054153
transform 1 0 6528 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1533
timestamp 1018054153
transform 1 0 6544 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1535
timestamp 1018054153
transform 1 0 6560 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1537
timestamp 1018054153
transform 1 0 6576 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1539
timestamp 1018054153
transform 1 0 6592 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1541
timestamp 1018054153
transform 1 0 6608 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1543
timestamp 1018054153
transform 1 0 6624 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1545
timestamp 1018054153
transform 1 0 6640 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1547
timestamp 1018054153
transform 1 0 6656 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1549
timestamp 1018054153
transform 1 0 6672 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1551
timestamp 1018054153
transform 1 0 6688 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1553
timestamp 1018054153
transform 1 0 6704 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1555
timestamp 1018054153
transform 1 0 6720 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1557
timestamp 1018054153
transform 1 0 6736 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1559
timestamp 1018054153
transform 1 0 6752 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1561
timestamp 1018054153
transform 1 0 6768 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1563
timestamp 1018054153
transform 1 0 6784 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1565
timestamp 1018054153
transform 1 0 6800 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1567
timestamp 1018054153
transform 1 0 6816 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1569
timestamp 1018054153
transform 1 0 6832 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1571
timestamp 1018054153
transform 1 0 6848 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1573
timestamp 1018054153
transform 1 0 6864 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1575
timestamp 1018054153
transform 1 0 6880 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1577
timestamp 1018054153
transform 1 0 6896 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1579
timestamp 1018054153
transform 1 0 6912 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1581
timestamp 1018054153
transform 1 0 6928 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1583
timestamp 1018054153
transform 1 0 6944 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1585
timestamp 1018054153
transform 1 0 6960 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1587
timestamp 1018054153
transform 1 0 6976 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1589
timestamp 1018054153
transform 1 0 6992 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1591
timestamp 1018054153
transform 1 0 7008 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1593
timestamp 1018054153
transform 1 0 7024 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1595
timestamp 1018054153
transform 1 0 7040 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1597
timestamp 1018054153
transform 1 0 7056 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1599
timestamp 1018054153
transform 1 0 7072 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1601
timestamp 1018054153
transform 1 0 7088 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1603
timestamp 1018054153
transform 1 0 7104 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1605
timestamp 1018054153
transform 1 0 7120 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1607
timestamp 1018054153
transform 1 0 7136 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1609
timestamp 1018054153
transform 1 0 7152 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1611
timestamp 1018054153
transform 1 0 7168 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1613
timestamp 1018054153
transform 1 0 7184 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1615
timestamp 1018054153
transform 1 0 7200 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1617
timestamp 1018054153
transform 1 0 7216 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1619
timestamp 1018054153
transform 1 0 7232 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1621
timestamp 1018054153
transform 1 0 7248 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1623
timestamp 1018054153
transform 1 0 7264 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1625
timestamp 1018054153
transform 1 0 7280 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1627
timestamp 1018054153
transform 1 0 7296 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1629
timestamp 1018054153
transform 1 0 7312 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1631
timestamp 1018054153
transform 1 0 7328 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1633
timestamp 1018054153
transform 1 0 7344 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1635
timestamp 1018054153
transform 1 0 7360 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1637
timestamp 1018054153
transform 1 0 7376 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1639
timestamp 1018054153
transform 1 0 7392 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1641
timestamp 1018054153
transform 1 0 7408 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1643
timestamp 1018054153
transform 1 0 7424 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1645
timestamp 1018054153
transform 1 0 7440 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1647
timestamp 1018054153
transform 1 0 7456 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1649
timestamp 1018054153
transform 1 0 7472 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1651
timestamp 1018054153
transform 1 0 7488 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1653
timestamp 1018054153
transform 1 0 7504 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1655
timestamp 1018054153
transform 1 0 7520 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1657
timestamp 1018054153
transform 1 0 7536 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1659
timestamp 1018054153
transform 1 0 7552 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1661
timestamp 1018054153
transform 1 0 7568 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1663
timestamp 1018054153
transform 1 0 7584 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1665
timestamp 1018054153
transform 1 0 7600 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1667
timestamp 1018054153
transform 1 0 7616 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1669
timestamp 1018054153
transform 1 0 7632 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1671
timestamp 1018054153
transform 1 0 7648 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1673
timestamp 1018054153
transform 1 0 7664 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1675
timestamp 1018054153
transform 1 0 7680 0 -1 6880
box -16 -6 32 210
use FILL  FILL_1677
timestamp 1018054153
transform 1 0 7696 0 -1 6880
box -16 -6 32 210
use PADVDD  PADVDD_0
timestamp 1084294447
transform 0 1 8000 -1 0 7400
box -6 -6 606 2000
use mult_pad_VIA1  mult_pad_VIA1_7
timestamp 1542725905
transform 1 0 7788 0 1 6680
box -48 -6 48 6
use FILL  FILL_1679
timestamp 1018054153
transform 1 0 7712 0 -1 6880
box -16 -6 32 210
use M2_M1  M2_M1_30
timestamp 1542725905
transform 1 0 3864 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_41
timestamp 1542725905
transform 1 0 3960 0 1 6530
box -4 -4 4 4
use M3_M2  M3_M2_5
timestamp 1542725905
transform 1 0 3960 0 1 6510
box -6 -6 6 6
use M3_M2  M3_M2_6
timestamp 1542725905
transform 1 0 4104 0 1 6510
box -6 -6 6 6
use M2_M1  M2_M1_24
timestamp 1542725905
transform 1 0 4344 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_31
timestamp 1542725905
transform 1 0 4344 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_19
timestamp 1542725905
transform 1 0 4392 0 1 6590
box -4 -4 4 4
use M2_M1  M2_M1_25
timestamp 1542725905
transform 1 0 4776 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_32
timestamp 1542725905
transform 1 0 4792 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_20
timestamp 1542725905
transform 1 0 4856 0 1 6590
box -4 -4 4 4
use M2_M1  M2_M1_26
timestamp 1542725905
transform 1 0 4824 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_27
timestamp 1542725905
transform 1 0 4856 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_33
timestamp 1542725905
transform 1 0 4856 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_21
timestamp 1542725905
transform 1 0 5080 0 1 6590
box -4 -4 4 4
use M2_M1  M2_M1_28
timestamp 1542725905
transform 1 0 5160 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_34
timestamp 1542725905
transform 1 0 5448 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_35
timestamp 1542725905
transform 1 0 5464 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_42
timestamp 1542725905
transform 1 0 5480 0 1 6530
box -4 -4 4 4
use M3_M2  M3_M2_7
timestamp 1542725905
transform 1 0 5496 0 1 6510
box -6 -6 6 6
use M2_M1  M2_M1_22
timestamp 1542725905
transform 1 0 5560 0 1 6590
box -4 -4 4 4
use M2_M1  M2_M1_36
timestamp 1542725905
transform 1 0 5704 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_37
timestamp 1542725905
transform 1 0 5768 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_38
timestamp 1542725905
transform 1 0 5960 0 1 6550
box -4 -4 4 4
use M2_M1  M2_M1_29
timestamp 1542725905
transform 1 0 6008 0 1 6570
box -4 -4 4 4
use M2_M1  M2_M1_23
timestamp 1542725905
transform 1 0 6280 0 1 6590
box -4 -4 4 4
use M2_M1  M2_M1_39
timestamp 1542725905
transform 1 0 6328 0 1 6550
box -4 -4 4 4
use M3_M2  M3_M2_4
timestamp 1542725905
transform 1 0 6328 0 1 6530
box -6 -6 6 6
use M2_M1  M2_M1_40
timestamp 1542725905
transform 1 0 6728 0 1 6550
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_8
timestamp 1542725905
transform 1 0 2092 0 1 6480
box -48 -6 48 6
use FILL  FILL_1680
timestamp 1018054153
transform 1 0 2272 0 1 6480
box -16 -6 32 210
use FILL  FILL_1682
timestamp 1018054153
transform 1 0 2288 0 1 6480
box -16 -6 32 210
use FILL  FILL_1684
timestamp 1018054153
transform 1 0 2304 0 1 6480
box -16 -6 32 210
use FILL  FILL_1686
timestamp 1018054153
transform 1 0 2320 0 1 6480
box -16 -6 32 210
use FILL  FILL_1688
timestamp 1018054153
transform 1 0 2336 0 1 6480
box -16 -6 32 210
use FILL  FILL_1690
timestamp 1018054153
transform 1 0 2352 0 1 6480
box -16 -6 32 210
use FILL  FILL_1692
timestamp 1018054153
transform 1 0 2368 0 1 6480
box -16 -6 32 210
use FILL  FILL_1694
timestamp 1018054153
transform 1 0 2384 0 1 6480
box -16 -6 32 210
use FILL  FILL_1696
timestamp 1018054153
transform 1 0 2400 0 1 6480
box -16 -6 32 210
use FILL  FILL_1698
timestamp 1018054153
transform 1 0 2416 0 1 6480
box -16 -6 32 210
use FILL  FILL_1700
timestamp 1018054153
transform 1 0 2432 0 1 6480
box -16 -6 32 210
use FILL  FILL_1702
timestamp 1018054153
transform 1 0 2448 0 1 6480
box -16 -6 32 210
use FILL  FILL_1704
timestamp 1018054153
transform 1 0 2464 0 1 6480
box -16 -6 32 210
use FILL  FILL_1706
timestamp 1018054153
transform 1 0 2480 0 1 6480
box -16 -6 32 210
use FILL  FILL_1708
timestamp 1018054153
transform 1 0 2496 0 1 6480
box -16 -6 32 210
use FILL  FILL_1710
timestamp 1018054153
transform 1 0 2512 0 1 6480
box -16 -6 32 210
use FILL  FILL_1712
timestamp 1018054153
transform 1 0 2528 0 1 6480
box -16 -6 32 210
use FILL  FILL_1714
timestamp 1018054153
transform 1 0 2544 0 1 6480
box -16 -6 32 210
use FILL  FILL_1716
timestamp 1018054153
transform 1 0 2560 0 1 6480
box -16 -6 32 210
use FILL  FILL_1718
timestamp 1018054153
transform 1 0 2576 0 1 6480
box -16 -6 32 210
use FILL  FILL_1720
timestamp 1018054153
transform 1 0 2592 0 1 6480
box -16 -6 32 210
use FILL  FILL_1722
timestamp 1018054153
transform 1 0 2608 0 1 6480
box -16 -6 32 210
use FILL  FILL_1724
timestamp 1018054153
transform 1 0 2624 0 1 6480
box -16 -6 32 210
use FILL  FILL_1726
timestamp 1018054153
transform 1 0 2640 0 1 6480
box -16 -6 32 210
use FILL  FILL_1728
timestamp 1018054153
transform 1 0 2656 0 1 6480
box -16 -6 32 210
use FILL  FILL_1730
timestamp 1018054153
transform 1 0 2672 0 1 6480
box -16 -6 32 210
use FILL  FILL_1732
timestamp 1018054153
transform 1 0 2688 0 1 6480
box -16 -6 32 210
use FILL  FILL_1734
timestamp 1018054153
transform 1 0 2704 0 1 6480
box -16 -6 32 210
use FILL  FILL_1736
timestamp 1018054153
transform 1 0 2720 0 1 6480
box -16 -6 32 210
use FILL  FILL_1738
timestamp 1018054153
transform 1 0 2736 0 1 6480
box -16 -6 32 210
use FILL  FILL_1740
timestamp 1018054153
transform 1 0 2752 0 1 6480
box -16 -6 32 210
use FILL  FILL_1742
timestamp 1018054153
transform 1 0 2768 0 1 6480
box -16 -6 32 210
use FILL  FILL_1744
timestamp 1018054153
transform 1 0 2784 0 1 6480
box -16 -6 32 210
use FILL  FILL_1746
timestamp 1018054153
transform 1 0 2800 0 1 6480
box -16 -6 32 210
use FILL  FILL_1748
timestamp 1018054153
transform 1 0 2816 0 1 6480
box -16 -6 32 210
use FILL  FILL_1750
timestamp 1018054153
transform 1 0 2832 0 1 6480
box -16 -6 32 210
use FILL  FILL_1752
timestamp 1018054153
transform 1 0 2848 0 1 6480
box -16 -6 32 210
use FILL  FILL_1754
timestamp 1018054153
transform 1 0 2864 0 1 6480
box -16 -6 32 210
use FILL  FILL_1756
timestamp 1018054153
transform 1 0 2880 0 1 6480
box -16 -6 32 210
use FILL  FILL_1758
timestamp 1018054153
transform 1 0 2896 0 1 6480
box -16 -6 32 210
use FILL  FILL_1760
timestamp 1018054153
transform 1 0 2912 0 1 6480
box -16 -6 32 210
use FILL  FILL_1762
timestamp 1018054153
transform 1 0 2928 0 1 6480
box -16 -6 32 210
use FILL  FILL_1764
timestamp 1018054153
transform 1 0 2944 0 1 6480
box -16 -6 32 210
use FILL  FILL_1766
timestamp 1018054153
transform 1 0 2960 0 1 6480
box -16 -6 32 210
use FILL  FILL_1768
timestamp 1018054153
transform 1 0 2976 0 1 6480
box -16 -6 32 210
use FILL  FILL_1770
timestamp 1018054153
transform 1 0 2992 0 1 6480
box -16 -6 32 210
use FILL  FILL_1772
timestamp 1018054153
transform 1 0 3008 0 1 6480
box -16 -6 32 210
use FILL  FILL_1774
timestamp 1018054153
transform 1 0 3024 0 1 6480
box -16 -6 32 210
use FILL  FILL_1776
timestamp 1018054153
transform 1 0 3040 0 1 6480
box -16 -6 32 210
use FILL  FILL_1778
timestamp 1018054153
transform 1 0 3056 0 1 6480
box -16 -6 32 210
use FILL  FILL_1780
timestamp 1018054153
transform 1 0 3072 0 1 6480
box -16 -6 32 210
use FILL  FILL_1782
timestamp 1018054153
transform 1 0 3088 0 1 6480
box -16 -6 32 210
use FILL  FILL_1784
timestamp 1018054153
transform 1 0 3104 0 1 6480
box -16 -6 32 210
use FILL  FILL_1786
timestamp 1018054153
transform 1 0 3120 0 1 6480
box -16 -6 32 210
use FILL  FILL_1788
timestamp 1018054153
transform 1 0 3136 0 1 6480
box -16 -6 32 210
use FILL  FILL_1790
timestamp 1018054153
transform 1 0 3152 0 1 6480
box -16 -6 32 210
use FILL  FILL_1792
timestamp 1018054153
transform 1 0 3168 0 1 6480
box -16 -6 32 210
use FILL  FILL_1794
timestamp 1018054153
transform 1 0 3184 0 1 6480
box -16 -6 32 210
use FILL  FILL_1796
timestamp 1018054153
transform 1 0 3200 0 1 6480
box -16 -6 32 210
use FILL  FILL_1798
timestamp 1018054153
transform 1 0 3216 0 1 6480
box -16 -6 32 210
use FILL  FILL_1800
timestamp 1018054153
transform 1 0 3232 0 1 6480
box -16 -6 32 210
use FILL  FILL_1802
timestamp 1018054153
transform 1 0 3248 0 1 6480
box -16 -6 32 210
use FILL  FILL_1804
timestamp 1018054153
transform 1 0 3264 0 1 6480
box -16 -6 32 210
use FILL  FILL_1806
timestamp 1018054153
transform 1 0 3280 0 1 6480
box -16 -6 32 210
use FILL  FILL_1808
timestamp 1018054153
transform 1 0 3296 0 1 6480
box -16 -6 32 210
use FILL  FILL_1810
timestamp 1018054153
transform 1 0 3312 0 1 6480
box -16 -6 32 210
use FILL  FILL_1812
timestamp 1018054153
transform 1 0 3328 0 1 6480
box -16 -6 32 210
use FILL  FILL_1814
timestamp 1018054153
transform 1 0 3344 0 1 6480
box -16 -6 32 210
use FILL  FILL_1816
timestamp 1018054153
transform 1 0 3360 0 1 6480
box -16 -6 32 210
use FILL  FILL_1818
timestamp 1018054153
transform 1 0 3376 0 1 6480
box -16 -6 32 210
use FILL  FILL_1820
timestamp 1018054153
transform 1 0 3392 0 1 6480
box -16 -6 32 210
use FILL  FILL_1822
timestamp 1018054153
transform 1 0 3408 0 1 6480
box -16 -6 32 210
use FILL  FILL_1824
timestamp 1018054153
transform 1 0 3424 0 1 6480
box -16 -6 32 210
use FILL  FILL_1826
timestamp 1018054153
transform 1 0 3440 0 1 6480
box -16 -6 32 210
use FILL  FILL_1828
timestamp 1018054153
transform 1 0 3456 0 1 6480
box -16 -6 32 210
use FILL  FILL_1830
timestamp 1018054153
transform 1 0 3472 0 1 6480
box -16 -6 32 210
use FILL  FILL_1832
timestamp 1018054153
transform 1 0 3488 0 1 6480
box -16 -6 32 210
use FILL  FILL_1834
timestamp 1018054153
transform 1 0 3504 0 1 6480
box -16 -6 32 210
use FILL  FILL_1836
timestamp 1018054153
transform 1 0 3520 0 1 6480
box -16 -6 32 210
use FILL  FILL_1838
timestamp 1018054153
transform 1 0 3536 0 1 6480
box -16 -6 32 210
use FILL  FILL_1840
timestamp 1018054153
transform 1 0 3552 0 1 6480
box -16 -6 32 210
use FILL  FILL_1842
timestamp 1018054153
transform 1 0 3568 0 1 6480
box -16 -6 32 210
use FILL  FILL_1844
timestamp 1018054153
transform 1 0 3584 0 1 6480
box -16 -6 32 210
use FILL  FILL_1846
timestamp 1018054153
transform 1 0 3600 0 1 6480
box -16 -6 32 210
use FILL  FILL_1848
timestamp 1018054153
transform 1 0 3616 0 1 6480
box -16 -6 32 210
use FILL  FILL_1850
timestamp 1018054153
transform 1 0 3632 0 1 6480
box -16 -6 32 210
use FILL  FILL_1852
timestamp 1018054153
transform 1 0 3648 0 1 6480
box -16 -6 32 210
use FILL  FILL_1854
timestamp 1018054153
transform 1 0 3664 0 1 6480
box -16 -6 32 210
use FILL  FILL_1856
timestamp 1018054153
transform 1 0 3680 0 1 6480
box -16 -6 32 210
use FILL  FILL_1858
timestamp 1018054153
transform 1 0 3696 0 1 6480
box -16 -6 32 210
use FILL  FILL_1860
timestamp 1018054153
transform 1 0 3712 0 1 6480
box -16 -6 32 210
use FILL  FILL_1862
timestamp 1018054153
transform 1 0 3728 0 1 6480
box -16 -6 32 210
use FILL  FILL_1864
timestamp 1018054153
transform 1 0 3744 0 1 6480
box -16 -6 32 210
use FILL  FILL_1866
timestamp 1018054153
transform 1 0 3760 0 1 6480
box -16 -6 32 210
use FILL  FILL_1868
timestamp 1018054153
transform 1 0 3776 0 1 6480
box -16 -6 32 210
use FILL  FILL_1870
timestamp 1018054153
transform 1 0 3792 0 1 6480
box -16 -6 32 210
use FILL  FILL_1872
timestamp 1018054153
transform 1 0 3808 0 1 6480
box -16 -6 32 210
use FILL  FILL_1873
timestamp 1018054153
transform 1 0 3824 0 1 6480
box -16 -6 32 210
use FILL  FILL_1874
timestamp 1018054153
transform 1 0 3840 0 1 6480
box -16 -6 32 210
use FILL  FILL_1875
timestamp 1018054153
transform 1 0 3856 0 1 6480
box -16 -6 32 210
use FILL  FILL_1877
timestamp 1018054153
transform 1 0 3872 0 1 6480
box -16 -6 32 210
use FILL  FILL_1879
timestamp 1018054153
transform 1 0 3888 0 1 6480
box -16 -6 32 210
use FILL  FILL_1881
timestamp 1018054153
transform 1 0 3904 0 1 6480
box -16 -6 32 210
use FILL  FILL_1883
timestamp 1018054153
transform 1 0 3920 0 1 6480
box -16 -6 32 210
use FILL  FILL_1885
timestamp 1018054153
transform 1 0 3936 0 1 6480
box -16 -6 32 210
use INVX1  INVX1_2
timestamp 1053022145
transform 1 0 3952 0 1 6480
box -18 -6 52 210
use FILL  FILL_1887
timestamp 1018054153
transform 1 0 3984 0 1 6480
box -16 -6 32 210
use FILL  FILL_1891
timestamp 1018054153
transform 1 0 4000 0 1 6480
box -16 -6 32 210
use FILL  FILL_1893
timestamp 1018054153
transform 1 0 4016 0 1 6480
box -16 -6 32 210
use FILL  FILL_1895
timestamp 1018054153
transform 1 0 4032 0 1 6480
box -16 -6 32 210
use FILL  FILL_1897
timestamp 1018054153
transform 1 0 4048 0 1 6480
box -16 -6 32 210
use FILL  FILL_1899
timestamp 1018054153
transform 1 0 4064 0 1 6480
box -16 -6 32 210
use FILL  FILL_1901
timestamp 1018054153
transform 1 0 4080 0 1 6480
box -16 -6 32 210
use FILL  FILL_1903
timestamp 1018054153
transform 1 0 4096 0 1 6480
box -16 -6 32 210
use FILL  FILL_1905
timestamp 1018054153
transform 1 0 4112 0 1 6480
box -16 -6 32 210
use FILL  FILL_1907
timestamp 1018054153
transform 1 0 4128 0 1 6480
box -16 -6 32 210
use FILL  FILL_1909
timestamp 1018054153
transform 1 0 4144 0 1 6480
box -16 -6 32 210
use FILL  FILL_1911
timestamp 1018054153
transform 1 0 4160 0 1 6480
box -16 -6 32 210
use FILL  FILL_1913
timestamp 1018054153
transform 1 0 4176 0 1 6480
box -16 -6 32 210
use FILL  FILL_1915
timestamp 1018054153
transform 1 0 4192 0 1 6480
box -16 -6 32 210
use FILL  FILL_1917
timestamp 1018054153
transform 1 0 4208 0 1 6480
box -16 -6 32 210
use FILL  FILL_1919
timestamp 1018054153
transform 1 0 4224 0 1 6480
box -16 -6 32 210
use FILL  FILL_1921
timestamp 1018054153
transform 1 0 4240 0 1 6480
box -16 -6 32 210
use FILL  FILL_1923
timestamp 1018054153
transform 1 0 4256 0 1 6480
box -16 -6 32 210
use FILL  FILL_1925
timestamp 1018054153
transform 1 0 4272 0 1 6480
box -16 -6 32 210
use FILL  FILL_1927
timestamp 1018054153
transform 1 0 4288 0 1 6480
box -16 -6 32 210
use FILL  FILL_1929
timestamp 1018054153
transform 1 0 4304 0 1 6480
box -16 -6 32 210
use FILL  FILL_1931
timestamp 1018054153
transform 1 0 4320 0 1 6480
box -16 -6 32 210
use OAI21X1  OAI21X1_2
timestamp 1053722159
transform 1 0 4336 0 1 6480
box -16 -6 68 210
use FILL  FILL_1933
timestamp 1018054153
transform 1 0 4400 0 1 6480
box -16 -6 32 210
use FILL  FILL_1934
timestamp 1018054153
transform 1 0 4416 0 1 6480
box -16 -6 32 210
use FILL  FILL_1935
timestamp 1018054153
transform 1 0 4432 0 1 6480
box -16 -6 32 210
use FILL  FILL_1936
timestamp 1018054153
transform 1 0 4448 0 1 6480
box -16 -6 32 210
use FILL  FILL_1943
timestamp 1018054153
transform 1 0 4464 0 1 6480
box -16 -6 32 210
use FILL  FILL_1945
timestamp 1018054153
transform 1 0 4480 0 1 6480
box -16 -6 32 210
use FILL  FILL_1947
timestamp 1018054153
transform 1 0 4496 0 1 6480
box -16 -6 32 210
use FILL  FILL_1949
timestamp 1018054153
transform 1 0 4512 0 1 6480
box -16 -6 32 210
use FILL  FILL_1951
timestamp 1018054153
transform 1 0 4528 0 1 6480
box -16 -6 32 210
use FILL  FILL_1953
timestamp 1018054153
transform 1 0 4544 0 1 6480
box -16 -6 32 210
use FILL  FILL_1955
timestamp 1018054153
transform 1 0 4560 0 1 6480
box -16 -6 32 210
use FILL  FILL_1957
timestamp 1018054153
transform 1 0 4576 0 1 6480
box -16 -6 32 210
use FILL  FILL_1959
timestamp 1018054153
transform 1 0 4592 0 1 6480
box -16 -6 32 210
use FILL  FILL_1961
timestamp 1018054153
transform 1 0 4608 0 1 6480
box -16 -6 32 210
use FILL  FILL_1963
timestamp 1018054153
transform 1 0 4624 0 1 6480
box -16 -6 32 210
use FILL  FILL_1965
timestamp 1018054153
transform 1 0 4640 0 1 6480
box -16 -6 32 210
use FILL  FILL_1967
timestamp 1018054153
transform 1 0 4656 0 1 6480
box -16 -6 32 210
use FILL  FILL_1969
timestamp 1018054153
transform 1 0 4672 0 1 6480
box -16 -6 32 210
use FILL  FILL_1971
timestamp 1018054153
transform 1 0 4688 0 1 6480
box -16 -6 32 210
use FILL  FILL_1973
timestamp 1018054153
transform 1 0 4704 0 1 6480
box -16 -6 32 210
use FILL  FILL_1975
timestamp 1018054153
transform 1 0 4720 0 1 6480
box -16 -6 32 210
use FILL  FILL_1977
timestamp 1018054153
transform 1 0 4736 0 1 6480
box -16 -6 32 210
use FILL  FILL_1978
timestamp 1018054153
transform 1 0 4752 0 1 6480
box -16 -6 32 210
use FILL  FILL_1979
timestamp 1018054153
transform 1 0 4768 0 1 6480
box -16 -6 32 210
use FILL  FILL_1980
timestamp 1018054153
transform 1 0 4784 0 1 6480
box -16 -6 32 210
use OAI21X1  OAI21X1_3
timestamp 1053722159
transform 1 0 4800 0 1 6480
box -16 -6 68 210
use FILL  FILL_1981
timestamp 1018054153
transform 1 0 4864 0 1 6480
box -16 -6 32 210
use FILL  FILL_1988
timestamp 1018054153
transform 1 0 4880 0 1 6480
box -16 -6 32 210
use FILL  FILL_1990
timestamp 1018054153
transform 1 0 4896 0 1 6480
box -16 -6 32 210
use FILL  FILL_1992
timestamp 1018054153
transform 1 0 4912 0 1 6480
box -16 -6 32 210
use FILL  FILL_1994
timestamp 1018054153
transform 1 0 4928 0 1 6480
box -16 -6 32 210
use FILL  FILL_1996
timestamp 1018054153
transform 1 0 4944 0 1 6480
box -16 -6 32 210
use FILL  FILL_1998
timestamp 1018054153
transform 1 0 4960 0 1 6480
box -16 -6 32 210
use FILL  FILL_2000
timestamp 1018054153
transform 1 0 4976 0 1 6480
box -16 -6 32 210
use FILL  FILL_2002
timestamp 1018054153
transform 1 0 4992 0 1 6480
box -16 -6 32 210
use FILL  FILL_2004
timestamp 1018054153
transform 1 0 5008 0 1 6480
box -16 -6 32 210
use FILL  FILL_2006
timestamp 1018054153
transform 1 0 5024 0 1 6480
box -16 -6 32 210
use FILL  FILL_2008
timestamp 1018054153
transform 1 0 5040 0 1 6480
box -16 -6 32 210
use M3_M2  M3_M2_8
timestamp 1542725905
transform 1 0 5080 0 1 6490
box -6 -6 6 6
use FILL  FILL_2010
timestamp 1018054153
transform 1 0 5056 0 1 6480
box -16 -6 32 210
use FILL  FILL_2012
timestamp 1018054153
transform 1 0 5072 0 1 6480
box -16 -6 32 210
use FILL  FILL_2014
timestamp 1018054153
transform 1 0 5088 0 1 6480
box -16 -6 32 210
use FILL  FILL_2016
timestamp 1018054153
transform 1 0 5104 0 1 6480
box -16 -6 32 210
use FILL  FILL_2018
timestamp 1018054153
transform 1 0 5120 0 1 6480
box -16 -6 32 210
use FILL  FILL_2019
timestamp 1018054153
transform 1 0 5136 0 1 6480
box -16 -6 32 210
use FILL  FILL_2020
timestamp 1018054153
transform 1 0 5152 0 1 6480
box -16 -6 32 210
use FILL  FILL_2021
timestamp 1018054153
transform 1 0 5168 0 1 6480
box -16 -6 32 210
use FILL  FILL_2023
timestamp 1018054153
transform 1 0 5184 0 1 6480
box -16 -6 32 210
use NAND2X1  NAND2X1_3
timestamp 1053022145
transform -1 0 5248 0 1 6480
box -16 -6 64 210
use FILL  FILL_2024
timestamp 1018054153
transform 1 0 5248 0 1 6480
box -16 -6 32 210
use FILL  FILL_2030
timestamp 1018054153
transform 1 0 5264 0 1 6480
box -16 -6 32 210
use FILL  FILL_2032
timestamp 1018054153
transform 1 0 5280 0 1 6480
box -16 -6 32 210
use FILL  FILL_2034
timestamp 1018054153
transform 1 0 5296 0 1 6480
box -16 -6 32 210
use FILL  FILL_2036
timestamp 1018054153
transform 1 0 5312 0 1 6480
box -16 -6 32 210
use FILL  FILL_2038
timestamp 1018054153
transform 1 0 5328 0 1 6480
box -16 -6 32 210
use FILL  FILL_2040
timestamp 1018054153
transform 1 0 5344 0 1 6480
box -16 -6 32 210
use FILL  FILL_2042
timestamp 1018054153
transform 1 0 5360 0 1 6480
box -16 -6 32 210
use FILL  FILL_2044
timestamp 1018054153
transform 1 0 5376 0 1 6480
box -16 -6 32 210
use FILL  FILL_2046
timestamp 1018054153
transform 1 0 5392 0 1 6480
box -16 -6 32 210
use FILL  FILL_2048
timestamp 1018054153
transform 1 0 5408 0 1 6480
box -16 -6 32 210
use FILL  FILL_2050
timestamp 1018054153
transform 1 0 5424 0 1 6480
box -16 -6 32 210
use FILL  FILL_2051
timestamp 1018054153
transform 1 0 5440 0 1 6480
box -16 -6 32 210
use INVX1  INVX1_4
timestamp 1053022145
transform -1 0 5488 0 1 6480
box -18 -6 52 210
use FILL  FILL_2052
timestamp 1018054153
transform 1 0 5488 0 1 6480
box -16 -6 32 210
use FILL  FILL_2054
timestamp 1018054153
transform 1 0 5504 0 1 6480
box -16 -6 32 210
use FILL  FILL_2056
timestamp 1018054153
transform 1 0 5520 0 1 6480
box -16 -6 32 210
use FILL  FILL_2058
timestamp 1018054153
transform 1 0 5536 0 1 6480
box -16 -6 32 210
use FILL  FILL_2060
timestamp 1018054153
transform 1 0 5552 0 1 6480
box -16 -6 32 210
use FILL  FILL_2062
timestamp 1018054153
transform 1 0 5568 0 1 6480
box -16 -6 32 210
use FILL  FILL_2064
timestamp 1018054153
transform 1 0 5584 0 1 6480
box -16 -6 32 210
use FILL  FILL_2066
timestamp 1018054153
transform 1 0 5600 0 1 6480
box -16 -6 32 210
use FILL  FILL_2068
timestamp 1018054153
transform 1 0 5616 0 1 6480
box -16 -6 32 210
use FILL  FILL_2070
timestamp 1018054153
transform 1 0 5632 0 1 6480
box -16 -6 32 210
use FILL  FILL_2072
timestamp 1018054153
transform 1 0 5648 0 1 6480
box -16 -6 32 210
use NAND2X1  NAND2X1_4
timestamp 1053022145
transform -1 0 5712 0 1 6480
box -16 -6 64 210
use FILL  FILL_2073
timestamp 1018054153
transform 1 0 5712 0 1 6480
box -16 -6 32 210
use FILL  FILL_2079
timestamp 1018054153
transform 1 0 5728 0 1 6480
box -16 -6 32 210
use FILL  FILL_2081
timestamp 1018054153
transform 1 0 5744 0 1 6480
box -16 -6 32 210
use FILL  FILL_2083
timestamp 1018054153
transform 1 0 5760 0 1 6480
box -16 -6 32 210
use FILL  FILL_2085
timestamp 1018054153
transform 1 0 5776 0 1 6480
box -16 -6 32 210
use FILL  FILL_2087
timestamp 1018054153
transform 1 0 5792 0 1 6480
box -16 -6 32 210
use FILL  FILL_2089
timestamp 1018054153
transform 1 0 5808 0 1 6480
box -16 -6 32 210
use FILL  FILL_2091
timestamp 1018054153
transform 1 0 5824 0 1 6480
box -16 -6 32 210
use FILL  FILL_2093
timestamp 1018054153
transform 1 0 5840 0 1 6480
box -16 -6 32 210
use FILL  FILL_2095
timestamp 1018054153
transform 1 0 5856 0 1 6480
box -16 -6 32 210
use FILL  FILL_2097
timestamp 1018054153
transform 1 0 5872 0 1 6480
box -16 -6 32 210
use OAI21X1  OAI21X1_5
timestamp 1053722159
transform -1 0 5952 0 1 6480
box -16 -6 68 210
use FILL  FILL_2098
timestamp 1018054153
transform 1 0 5952 0 1 6480
box -16 -6 32 210
use FILL  FILL_2099
timestamp 1018054153
transform 1 0 5968 0 1 6480
box -16 -6 32 210
use FILL  FILL_2100
timestamp 1018054153
transform 1 0 5984 0 1 6480
box -16 -6 32 210
use FILL  FILL_2105
timestamp 1018054153
transform 1 0 6000 0 1 6480
box -16 -6 32 210
use FILL  FILL_2107
timestamp 1018054153
transform 1 0 6016 0 1 6480
box -16 -6 32 210
use FILL  FILL_2109
timestamp 1018054153
transform 1 0 6032 0 1 6480
box -16 -6 32 210
use FILL  FILL_2111
timestamp 1018054153
transform 1 0 6048 0 1 6480
box -16 -6 32 210
use FILL  FILL_2113
timestamp 1018054153
transform 1 0 6064 0 1 6480
box -16 -6 32 210
use FILL  FILL_2115
timestamp 1018054153
transform 1 0 6080 0 1 6480
box -16 -6 32 210
use FILL  FILL_2117
timestamp 1018054153
transform 1 0 6096 0 1 6480
box -16 -6 32 210
use FILL  FILL_2119
timestamp 1018054153
transform 1 0 6112 0 1 6480
box -16 -6 32 210
use FILL  FILL_2121
timestamp 1018054153
transform 1 0 6128 0 1 6480
box -16 -6 32 210
use FILL  FILL_2123
timestamp 1018054153
transform 1 0 6144 0 1 6480
box -16 -6 32 210
use FILL  FILL_2125
timestamp 1018054153
transform 1 0 6160 0 1 6480
box -16 -6 32 210
use FILL  FILL_2127
timestamp 1018054153
transform 1 0 6176 0 1 6480
box -16 -6 32 210
use FILL  FILL_2129
timestamp 1018054153
transform 1 0 6192 0 1 6480
box -16 -6 32 210
use FILL  FILL_2131
timestamp 1018054153
transform 1 0 6208 0 1 6480
box -16 -6 32 210
use FILL  FILL_2133
timestamp 1018054153
transform 1 0 6224 0 1 6480
box -16 -6 32 210
use FILL  FILL_2135
timestamp 1018054153
transform 1 0 6240 0 1 6480
box -16 -6 32 210
use FILL  FILL_2137
timestamp 1018054153
transform 1 0 6256 0 1 6480
box -16 -6 32 210
use FILL  FILL_2139
timestamp 1018054153
transform 1 0 6272 0 1 6480
box -16 -6 32 210
use NAND2X1  NAND2X1_5
timestamp 1053022145
transform -1 0 6336 0 1 6480
box -16 -6 64 210
use FILL  FILL_2140
timestamp 1018054153
transform 1 0 6336 0 1 6480
box -16 -6 32 210
use FILL  FILL_2146
timestamp 1018054153
transform 1 0 6352 0 1 6480
box -16 -6 32 210
use FILL  FILL_2148
timestamp 1018054153
transform 1 0 6368 0 1 6480
box -16 -6 32 210
use FILL  FILL_2150
timestamp 1018054153
transform 1 0 6384 0 1 6480
box -16 -6 32 210
use FILL  FILL_2152
timestamp 1018054153
transform 1 0 6400 0 1 6480
box -16 -6 32 210
use FILL  FILL_2154
timestamp 1018054153
transform 1 0 6416 0 1 6480
box -16 -6 32 210
use FILL  FILL_2156
timestamp 1018054153
transform 1 0 6432 0 1 6480
box -16 -6 32 210
use FILL  FILL_2158
timestamp 1018054153
transform 1 0 6448 0 1 6480
box -16 -6 32 210
use FILL  FILL_2160
timestamp 1018054153
transform 1 0 6464 0 1 6480
box -16 -6 32 210
use FILL  FILL_2162
timestamp 1018054153
transform 1 0 6480 0 1 6480
box -16 -6 32 210
use FILL  FILL_2164
timestamp 1018054153
transform 1 0 6496 0 1 6480
box -16 -6 32 210
use FILL  FILL_2166
timestamp 1018054153
transform 1 0 6512 0 1 6480
box -16 -6 32 210
use FILL  FILL_2168
timestamp 1018054153
transform 1 0 6528 0 1 6480
box -16 -6 32 210
use FILL  FILL_2170
timestamp 1018054153
transform 1 0 6544 0 1 6480
box -16 -6 32 210
use FILL  FILL_2172
timestamp 1018054153
transform 1 0 6560 0 1 6480
box -16 -6 32 210
use FILL  FILL_2174
timestamp 1018054153
transform 1 0 6576 0 1 6480
box -16 -6 32 210
use FILL  FILL_2176
timestamp 1018054153
transform 1 0 6592 0 1 6480
box -16 -6 32 210
use FILL  FILL_2178
timestamp 1018054153
transform 1 0 6608 0 1 6480
box -16 -6 32 210
use FILL  FILL_2180
timestamp 1018054153
transform 1 0 6624 0 1 6480
box -16 -6 32 210
use FILL  FILL_2182
timestamp 1018054153
transform 1 0 6640 0 1 6480
box -16 -6 32 210
use FILL  FILL_2184
timestamp 1018054153
transform 1 0 6656 0 1 6480
box -16 -6 32 210
use FILL  FILL_2186
timestamp 1018054153
transform 1 0 6672 0 1 6480
box -16 -6 32 210
use FILL  FILL_2188
timestamp 1018054153
transform 1 0 6688 0 1 6480
box -16 -6 32 210
use FILL  FILL_2190
timestamp 1018054153
transform 1 0 6704 0 1 6480
box -16 -6 32 210
use FILL  FILL_2192
timestamp 1018054153
transform 1 0 6720 0 1 6480
box -16 -6 32 210
use FILL  FILL_2194
timestamp 1018054153
transform 1 0 6736 0 1 6480
box -16 -6 32 210
use FILL  FILL_2196
timestamp 1018054153
transform 1 0 6752 0 1 6480
box -16 -6 32 210
use FILL  FILL_2198
timestamp 1018054153
transform 1 0 6768 0 1 6480
box -16 -6 32 210
use FILL  FILL_2200
timestamp 1018054153
transform 1 0 6784 0 1 6480
box -16 -6 32 210
use FILL  FILL_2202
timestamp 1018054153
transform 1 0 6800 0 1 6480
box -16 -6 32 210
use FILL  FILL_2204
timestamp 1018054153
transform 1 0 6816 0 1 6480
box -16 -6 32 210
use FILL  FILL_2206
timestamp 1018054153
transform 1 0 6832 0 1 6480
box -16 -6 32 210
use FILL  FILL_2208
timestamp 1018054153
transform 1 0 6848 0 1 6480
box -16 -6 32 210
use FILL  FILL_2210
timestamp 1018054153
transform 1 0 6864 0 1 6480
box -16 -6 32 210
use FILL  FILL_2212
timestamp 1018054153
transform 1 0 6880 0 1 6480
box -16 -6 32 210
use FILL  FILL_2214
timestamp 1018054153
transform 1 0 6896 0 1 6480
box -16 -6 32 210
use FILL  FILL_2216
timestamp 1018054153
transform 1 0 6912 0 1 6480
box -16 -6 32 210
use FILL  FILL_2218
timestamp 1018054153
transform 1 0 6928 0 1 6480
box -16 -6 32 210
use FILL  FILL_2220
timestamp 1018054153
transform 1 0 6944 0 1 6480
box -16 -6 32 210
use FILL  FILL_2222
timestamp 1018054153
transform 1 0 6960 0 1 6480
box -16 -6 32 210
use FILL  FILL_2224
timestamp 1018054153
transform 1 0 6976 0 1 6480
box -16 -6 32 210
use FILL  FILL_2226
timestamp 1018054153
transform 1 0 6992 0 1 6480
box -16 -6 32 210
use FILL  FILL_2228
timestamp 1018054153
transform 1 0 7008 0 1 6480
box -16 -6 32 210
use FILL  FILL_2230
timestamp 1018054153
transform 1 0 7024 0 1 6480
box -16 -6 32 210
use FILL  FILL_2232
timestamp 1018054153
transform 1 0 7040 0 1 6480
box -16 -6 32 210
use FILL  FILL_2234
timestamp 1018054153
transform 1 0 7056 0 1 6480
box -16 -6 32 210
use FILL  FILL_2236
timestamp 1018054153
transform 1 0 7072 0 1 6480
box -16 -6 32 210
use FILL  FILL_2238
timestamp 1018054153
transform 1 0 7088 0 1 6480
box -16 -6 32 210
use FILL  FILL_2240
timestamp 1018054153
transform 1 0 7104 0 1 6480
box -16 -6 32 210
use FILL  FILL_2242
timestamp 1018054153
transform 1 0 7120 0 1 6480
box -16 -6 32 210
use FILL  FILL_2244
timestamp 1018054153
transform 1 0 7136 0 1 6480
box -16 -6 32 210
use FILL  FILL_2246
timestamp 1018054153
transform 1 0 7152 0 1 6480
box -16 -6 32 210
use FILL  FILL_2248
timestamp 1018054153
transform 1 0 7168 0 1 6480
box -16 -6 32 210
use FILL  FILL_2250
timestamp 1018054153
transform 1 0 7184 0 1 6480
box -16 -6 32 210
use FILL  FILL_2252
timestamp 1018054153
transform 1 0 7200 0 1 6480
box -16 -6 32 210
use FILL  FILL_2254
timestamp 1018054153
transform 1 0 7216 0 1 6480
box -16 -6 32 210
use FILL  FILL_2256
timestamp 1018054153
transform 1 0 7232 0 1 6480
box -16 -6 32 210
use FILL  FILL_2258
timestamp 1018054153
transform 1 0 7248 0 1 6480
box -16 -6 32 210
use FILL  FILL_2260
timestamp 1018054153
transform 1 0 7264 0 1 6480
box -16 -6 32 210
use FILL  FILL_2262
timestamp 1018054153
transform 1 0 7280 0 1 6480
box -16 -6 32 210
use FILL  FILL_2264
timestamp 1018054153
transform 1 0 7296 0 1 6480
box -16 -6 32 210
use FILL  FILL_2266
timestamp 1018054153
transform 1 0 7312 0 1 6480
box -16 -6 32 210
use FILL  FILL_2268
timestamp 1018054153
transform 1 0 7328 0 1 6480
box -16 -6 32 210
use FILL  FILL_2270
timestamp 1018054153
transform 1 0 7344 0 1 6480
box -16 -6 32 210
use FILL  FILL_2272
timestamp 1018054153
transform 1 0 7360 0 1 6480
box -16 -6 32 210
use FILL  FILL_2274
timestamp 1018054153
transform 1 0 7376 0 1 6480
box -16 -6 32 210
use FILL  FILL_2276
timestamp 1018054153
transform 1 0 7392 0 1 6480
box -16 -6 32 210
use FILL  FILL_2278
timestamp 1018054153
transform 1 0 7408 0 1 6480
box -16 -6 32 210
use FILL  FILL_2280
timestamp 1018054153
transform 1 0 7424 0 1 6480
box -16 -6 32 210
use FILL  FILL_2282
timestamp 1018054153
transform 1 0 7440 0 1 6480
box -16 -6 32 210
use FILL  FILL_2284
timestamp 1018054153
transform 1 0 7456 0 1 6480
box -16 -6 32 210
use FILL  FILL_2286
timestamp 1018054153
transform 1 0 7472 0 1 6480
box -16 -6 32 210
use FILL  FILL_2288
timestamp 1018054153
transform 1 0 7488 0 1 6480
box -16 -6 32 210
use FILL  FILL_2290
timestamp 1018054153
transform 1 0 7504 0 1 6480
box -16 -6 32 210
use FILL  FILL_2292
timestamp 1018054153
transform 1 0 7520 0 1 6480
box -16 -6 32 210
use FILL  FILL_2294
timestamp 1018054153
transform 1 0 7536 0 1 6480
box -16 -6 32 210
use FILL  FILL_2296
timestamp 1018054153
transform 1 0 7552 0 1 6480
box -16 -6 32 210
use FILL  FILL_2298
timestamp 1018054153
transform 1 0 7568 0 1 6480
box -16 -6 32 210
use FILL  FILL_2300
timestamp 1018054153
transform 1 0 7584 0 1 6480
box -16 -6 32 210
use FILL  FILL_2302
timestamp 1018054153
transform 1 0 7600 0 1 6480
box -16 -6 32 210
use FILL  FILL_2304
timestamp 1018054153
transform 1 0 7616 0 1 6480
box -16 -6 32 210
use FILL  FILL_2306
timestamp 1018054153
transform 1 0 7632 0 1 6480
box -16 -6 32 210
use FILL  FILL_2308
timestamp 1018054153
transform 1 0 7648 0 1 6480
box -16 -6 32 210
use FILL  FILL_2310
timestamp 1018054153
transform 1 0 7664 0 1 6480
box -16 -6 32 210
use FILL  FILL_2312
timestamp 1018054153
transform 1 0 7680 0 1 6480
box -16 -6 32 210
use FILL  FILL_2314
timestamp 1018054153
transform 1 0 7696 0 1 6480
box -16 -6 32 210
use FILL  FILL_2316
timestamp 1018054153
transform 1 0 7712 0 1 6480
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_9
timestamp 1542725905
transform 1 0 7908 0 1 6480
box -48 -6 48 6
use M2_M1  M2_M1_46
timestamp 1542725905
transform 1 0 3432 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_43
timestamp 1542725905
transform 1 0 3816 0 1 6430
box -4 -4 4 4
use M3_M2  M3_M2_9
timestamp 1542725905
transform 1 0 3832 0 1 6430
box -6 -6 6 6
use M2_M1  M2_M1_55
timestamp 1542725905
transform 1 0 3864 0 1 6390
box -4 -4 4 4
use M3_M2  M3_M2_10
timestamp 1542725905
transform 1 0 3928 0 1 6430
box -6 -6 6 6
use M2_M1  M2_M1_47
timestamp 1542725905
transform 1 0 3928 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_48
timestamp 1542725905
transform 1 0 4184 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_44
timestamp 1542725905
transform 1 0 4456 0 1 6430
box -4 -4 4 4
use M2_M1  M2_M1_56
timestamp 1542725905
transform 1 0 4440 0 1 6390
box -4 -4 4 4
use M2_M1  M2_M1_49
timestamp 1542725905
transform 1 0 4776 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_45
timestamp 1542725905
transform 1 0 4808 0 1 6430
box -4 -4 4 4
use M2_M1  M2_M1_50
timestamp 1542725905
transform 1 0 4856 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_51
timestamp 1542725905
transform 1 0 5064 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_60
timestamp 1542725905
transform 1 0 5160 0 1 6370
box -4 -4 4 4
use M2_M1  M2_M1_57
timestamp 1542725905
transform 1 0 5224 0 1 6390
box -4 -4 4 4
use M2_M1  M2_M1_52
timestamp 1542725905
transform 1 0 5400 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_58
timestamp 1542725905
transform 1 0 5432 0 1 6390
box -4 -4 4 4
use M2_M1  M2_M1_61
timestamp 1542725905
transform 1 0 5480 0 1 6370
box -4 -4 4 4
use M3_M2  M3_M2_11
timestamp 1542725905
transform 1 0 5624 0 1 6410
box -6 -6 6 6
use M2_M1  M2_M1_53
timestamp 1542725905
transform 1 0 5704 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_54
timestamp 1542725905
transform 1 0 5976 0 1 6410
box -4 -4 4 4
use M2_M1  M2_M1_59
timestamp 1542725905
transform 1 0 5960 0 1 6390
box -4 -4 4 4
use M3_M2  M3_M2_12
timestamp 1542725905
transform 1 0 6392 0 1 6410
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_10
timestamp 1542725905
transform 1 0 2212 0 1 6280
box -48 -6 48 6
use PADINC  PADINC_4
timestamp 1084294328
transform 0 -1 2000 1 0 6200
box -12 -6 606 2000
use M3_M2  M3_M2_23
timestamp 1542725905
transform 1 0 1998 0 1 6130
box -6 -6 6 6
use FILL  FILL_1681
timestamp 1018054153
transform 1 0 2272 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1683
timestamp 1018054153
transform 1 0 2288 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1685
timestamp 1018054153
transform 1 0 2304 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1687
timestamp 1018054153
transform 1 0 2320 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1689
timestamp 1018054153
transform 1 0 2336 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1691
timestamp 1018054153
transform 1 0 2352 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1693
timestamp 1018054153
transform 1 0 2368 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1695
timestamp 1018054153
transform 1 0 2384 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1697
timestamp 1018054153
transform 1 0 2400 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1699
timestamp 1018054153
transform 1 0 2416 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1701
timestamp 1018054153
transform 1 0 2432 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1703
timestamp 1018054153
transform 1 0 2448 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1705
timestamp 1018054153
transform 1 0 2464 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1707
timestamp 1018054153
transform 1 0 2480 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1709
timestamp 1018054153
transform 1 0 2496 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1711
timestamp 1018054153
transform 1 0 2512 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1713
timestamp 1018054153
transform 1 0 2528 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1715
timestamp 1018054153
transform 1 0 2544 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1717
timestamp 1018054153
transform 1 0 2560 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1719
timestamp 1018054153
transform 1 0 2576 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1721
timestamp 1018054153
transform 1 0 2592 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1723
timestamp 1018054153
transform 1 0 2608 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1725
timestamp 1018054153
transform 1 0 2624 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1727
timestamp 1018054153
transform 1 0 2640 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1729
timestamp 1018054153
transform 1 0 2656 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1731
timestamp 1018054153
transform 1 0 2672 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1733
timestamp 1018054153
transform 1 0 2688 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1735
timestamp 1018054153
transform 1 0 2704 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1737
timestamp 1018054153
transform 1 0 2720 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1739
timestamp 1018054153
transform 1 0 2736 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1741
timestamp 1018054153
transform 1 0 2752 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1743
timestamp 1018054153
transform 1 0 2768 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1745
timestamp 1018054153
transform 1 0 2784 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1747
timestamp 1018054153
transform 1 0 2800 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1749
timestamp 1018054153
transform 1 0 2816 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1751
timestamp 1018054153
transform 1 0 2832 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1753
timestamp 1018054153
transform 1 0 2848 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1755
timestamp 1018054153
transform 1 0 2864 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1757
timestamp 1018054153
transform 1 0 2880 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1759
timestamp 1018054153
transform 1 0 2896 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1761
timestamp 1018054153
transform 1 0 2912 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1763
timestamp 1018054153
transform 1 0 2928 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1765
timestamp 1018054153
transform 1 0 2944 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1767
timestamp 1018054153
transform 1 0 2960 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1769
timestamp 1018054153
transform 1 0 2976 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1771
timestamp 1018054153
transform 1 0 2992 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1773
timestamp 1018054153
transform 1 0 3008 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1775
timestamp 1018054153
transform 1 0 3024 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1777
timestamp 1018054153
transform 1 0 3040 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1779
timestamp 1018054153
transform 1 0 3056 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1781
timestamp 1018054153
transform 1 0 3072 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1783
timestamp 1018054153
transform 1 0 3088 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1785
timestamp 1018054153
transform 1 0 3104 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1787
timestamp 1018054153
transform 1 0 3120 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1789
timestamp 1018054153
transform 1 0 3136 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1791
timestamp 1018054153
transform 1 0 3152 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1793
timestamp 1018054153
transform 1 0 3168 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1795
timestamp 1018054153
transform 1 0 3184 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1797
timestamp 1018054153
transform 1 0 3200 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1799
timestamp 1018054153
transform 1 0 3216 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1801
timestamp 1018054153
transform 1 0 3232 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1803
timestamp 1018054153
transform 1 0 3248 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1805
timestamp 1018054153
transform 1 0 3264 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1807
timestamp 1018054153
transform 1 0 3280 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1809
timestamp 1018054153
transform 1 0 3296 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1811
timestamp 1018054153
transform 1 0 3312 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1813
timestamp 1018054153
transform 1 0 3328 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1815
timestamp 1018054153
transform 1 0 3344 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1817
timestamp 1018054153
transform 1 0 3360 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1819
timestamp 1018054153
transform 1 0 3376 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1821
timestamp 1018054153
transform 1 0 3392 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1823
timestamp 1018054153
transform 1 0 3408 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1825
timestamp 1018054153
transform 1 0 3424 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1827
timestamp 1018054153
transform 1 0 3440 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1829
timestamp 1018054153
transform 1 0 3456 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1831
timestamp 1018054153
transform 1 0 3472 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1833
timestamp 1018054153
transform 1 0 3488 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1835
timestamp 1018054153
transform 1 0 3504 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1837
timestamp 1018054153
transform 1 0 3520 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1839
timestamp 1018054153
transform 1 0 3536 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1841
timestamp 1018054153
transform 1 0 3552 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1843
timestamp 1018054153
transform 1 0 3568 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1845
timestamp 1018054153
transform 1 0 3584 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1847
timestamp 1018054153
transform 1 0 3600 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1849
timestamp 1018054153
transform 1 0 3616 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1851
timestamp 1018054153
transform 1 0 3632 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1853
timestamp 1018054153
transform 1 0 3648 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1855
timestamp 1018054153
transform 1 0 3664 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1857
timestamp 1018054153
transform 1 0 3680 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1859
timestamp 1018054153
transform 1 0 3696 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1861
timestamp 1018054153
transform 1 0 3712 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1863
timestamp 1018054153
transform 1 0 3728 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1865
timestamp 1018054153
transform 1 0 3744 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1867
timestamp 1018054153
transform 1 0 3760 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1869
timestamp 1018054153
transform 1 0 3776 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1871
timestamp 1018054153
transform 1 0 3792 0 -1 6480
box -16 -6 32 210
use NOR2X1  NOR2X1_0
timestamp 1053022145
transform 1 0 3808 0 -1 6480
box -16 -6 64 210
use FILL  FILL_1876
timestamp 1018054153
transform 1 0 3856 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1878
timestamp 1018054153
transform 1 0 3872 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1880
timestamp 1018054153
transform 1 0 3888 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1882
timestamp 1018054153
transform 1 0 3904 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1884
timestamp 1018054153
transform 1 0 3920 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1886
timestamp 1018054153
transform 1 0 3936 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1888
timestamp 1018054153
transform 1 0 3952 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1889
timestamp 1018054153
transform 1 0 3968 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1890
timestamp 1018054153
transform 1 0 3984 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1892
timestamp 1018054153
transform 1 0 4000 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1894
timestamp 1018054153
transform 1 0 4016 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1896
timestamp 1018054153
transform 1 0 4032 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1898
timestamp 1018054153
transform 1 0 4048 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1900
timestamp 1018054153
transform 1 0 4064 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1902
timestamp 1018054153
transform 1 0 4080 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1904
timestamp 1018054153
transform 1 0 4096 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1906
timestamp 1018054153
transform 1 0 4112 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1908
timestamp 1018054153
transform 1 0 4128 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1910
timestamp 1018054153
transform 1 0 4144 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1912
timestamp 1018054153
transform 1 0 4160 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1914
timestamp 1018054153
transform 1 0 4176 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1916
timestamp 1018054153
transform 1 0 4192 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1918
timestamp 1018054153
transform 1 0 4208 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1920
timestamp 1018054153
transform 1 0 4224 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1922
timestamp 1018054153
transform 1 0 4240 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1924
timestamp 1018054153
transform 1 0 4256 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1926
timestamp 1018054153
transform 1 0 4272 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1928
timestamp 1018054153
transform 1 0 4288 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1930
timestamp 1018054153
transform 1 0 4304 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1932
timestamp 1018054153
transform 1 0 4320 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1937
timestamp 1018054153
transform 1 0 4336 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1938
timestamp 1018054153
transform 1 0 4352 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1939
timestamp 1018054153
transform 1 0 4368 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1940
timestamp 1018054153
transform 1 0 4384 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1941
timestamp 1018054153
transform 1 0 4400 0 -1 6480
box -16 -6 32 210
use INVX1  INVX1_3
timestamp 1053022145
transform -1 0 4448 0 -1 6480
box -18 -6 52 210
use FILL  FILL_1942
timestamp 1018054153
transform 1 0 4448 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1944
timestamp 1018054153
transform 1 0 4464 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1946
timestamp 1018054153
transform 1 0 4480 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1948
timestamp 1018054153
transform 1 0 4496 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1950
timestamp 1018054153
transform 1 0 4512 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1952
timestamp 1018054153
transform 1 0 4528 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1954
timestamp 1018054153
transform 1 0 4544 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1956
timestamp 1018054153
transform 1 0 4560 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1958
timestamp 1018054153
transform 1 0 4576 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1960
timestamp 1018054153
transform 1 0 4592 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1962
timestamp 1018054153
transform 1 0 4608 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1964
timestamp 1018054153
transform 1 0 4624 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1966
timestamp 1018054153
transform 1 0 4640 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1968
timestamp 1018054153
transform 1 0 4656 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1970
timestamp 1018054153
transform 1 0 4672 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1972
timestamp 1018054153
transform 1 0 4688 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1974
timestamp 1018054153
transform 1 0 4704 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1976
timestamp 1018054153
transform 1 0 4720 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1982
timestamp 1018054153
transform 1 0 4736 0 -1 6480
box -16 -6 32 210
use NOR2X1  NOR2X1_1
timestamp 1053022145
transform -1 0 4800 0 -1 6480
box -16 -6 64 210
use FILL  FILL_1983
timestamp 1018054153
transform 1 0 4800 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1984
timestamp 1018054153
transform 1 0 4816 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1985
timestamp 1018054153
transform 1 0 4832 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1986
timestamp 1018054153
transform 1 0 4848 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1987
timestamp 1018054153
transform 1 0 4864 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1989
timestamp 1018054153
transform 1 0 4880 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1991
timestamp 1018054153
transform 1 0 4896 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1993
timestamp 1018054153
transform 1 0 4912 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1995
timestamp 1018054153
transform 1 0 4928 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1997
timestamp 1018054153
transform 1 0 4944 0 -1 6480
box -16 -6 32 210
use FILL  FILL_1999
timestamp 1018054153
transform 1 0 4960 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2001
timestamp 1018054153
transform 1 0 4976 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2003
timestamp 1018054153
transform 1 0 4992 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2005
timestamp 1018054153
transform 1 0 5008 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2007
timestamp 1018054153
transform 1 0 5024 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2009
timestamp 1018054153
transform 1 0 5040 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2011
timestamp 1018054153
transform 1 0 5056 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2013
timestamp 1018054153
transform 1 0 5072 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2015
timestamp 1018054153
transform 1 0 5088 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2017
timestamp 1018054153
transform 1 0 5104 0 -1 6480
box -16 -6 32 210
use NAND2X1  NAND2X1_2
timestamp 1053022145
transform 1 0 5120 0 -1 6480
box -16 -6 64 210
use FILL  FILL_2022
timestamp 1018054153
transform 1 0 5168 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2025
timestamp 1018054153
transform 1 0 5184 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2026
timestamp 1018054153
transform 1 0 5200 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2027
timestamp 1018054153
transform 1 0 5216 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2028
timestamp 1018054153
transform 1 0 5232 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2029
timestamp 1018054153
transform 1 0 5248 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2031
timestamp 1018054153
transform 1 0 5264 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2033
timestamp 1018054153
transform 1 0 5280 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2035
timestamp 1018054153
transform 1 0 5296 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2037
timestamp 1018054153
transform 1 0 5312 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2039
timestamp 1018054153
transform 1 0 5328 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2041
timestamp 1018054153
transform 1 0 5344 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2043
timestamp 1018054153
transform 1 0 5360 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2045
timestamp 1018054153
transform 1 0 5376 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2047
timestamp 1018054153
transform 1 0 5392 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2049
timestamp 1018054153
transform 1 0 5408 0 -1 6480
box -16 -6 32 210
use OAI21X1  OAI21X1_4
timestamp 1053722159
transform 1 0 5424 0 -1 6480
box -16 -6 68 210
use FILL  FILL_2053
timestamp 1018054153
transform 1 0 5488 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2055
timestamp 1018054153
transform 1 0 5504 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2057
timestamp 1018054153
transform 1 0 5520 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2059
timestamp 1018054153
transform 1 0 5536 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2061
timestamp 1018054153
transform 1 0 5552 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2063
timestamp 1018054153
transform 1 0 5568 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2065
timestamp 1018054153
transform 1 0 5584 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2067
timestamp 1018054153
transform 1 0 5600 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2069
timestamp 1018054153
transform 1 0 5616 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2071
timestamp 1018054153
transform 1 0 5632 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2074
timestamp 1018054153
transform 1 0 5648 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2075
timestamp 1018054153
transform 1 0 5664 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2076
timestamp 1018054153
transform 1 0 5680 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2077
timestamp 1018054153
transform 1 0 5696 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2078
timestamp 1018054153
transform 1 0 5712 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2080
timestamp 1018054153
transform 1 0 5728 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2082
timestamp 1018054153
transform 1 0 5744 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2084
timestamp 1018054153
transform 1 0 5760 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2086
timestamp 1018054153
transform 1 0 5776 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2088
timestamp 1018054153
transform 1 0 5792 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2090
timestamp 1018054153
transform 1 0 5808 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2092
timestamp 1018054153
transform 1 0 5824 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2094
timestamp 1018054153
transform 1 0 5840 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2096
timestamp 1018054153
transform 1 0 5856 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2101
timestamp 1018054153
transform 1 0 5872 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2102
timestamp 1018054153
transform 1 0 5888 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2103
timestamp 1018054153
transform 1 0 5904 0 -1 6480
box -16 -6 32 210
use OAI21X1  OAI21X1_6
timestamp 1053722159
transform -1 0 5984 0 -1 6480
box -16 -6 68 210
use FILL  FILL_2104
timestamp 1018054153
transform 1 0 5984 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2106
timestamp 1018054153
transform 1 0 6000 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2108
timestamp 1018054153
transform 1 0 6016 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2110
timestamp 1018054153
transform 1 0 6032 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2112
timestamp 1018054153
transform 1 0 6048 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2114
timestamp 1018054153
transform 1 0 6064 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2116
timestamp 1018054153
transform 1 0 6080 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2118
timestamp 1018054153
transform 1 0 6096 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2120
timestamp 1018054153
transform 1 0 6112 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2122
timestamp 1018054153
transform 1 0 6128 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2124
timestamp 1018054153
transform 1 0 6144 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2126
timestamp 1018054153
transform 1 0 6160 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2128
timestamp 1018054153
transform 1 0 6176 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2130
timestamp 1018054153
transform 1 0 6192 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2132
timestamp 1018054153
transform 1 0 6208 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2134
timestamp 1018054153
transform 1 0 6224 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2136
timestamp 1018054153
transform 1 0 6240 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2138
timestamp 1018054153
transform 1 0 6256 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2141
timestamp 1018054153
transform 1 0 6272 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2142
timestamp 1018054153
transform 1 0 6288 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2143
timestamp 1018054153
transform 1 0 6304 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2144
timestamp 1018054153
transform 1 0 6320 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2145
timestamp 1018054153
transform 1 0 6336 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2147
timestamp 1018054153
transform 1 0 6352 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2149
timestamp 1018054153
transform 1 0 6368 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2151
timestamp 1018054153
transform 1 0 6384 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2153
timestamp 1018054153
transform 1 0 6400 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2155
timestamp 1018054153
transform 1 0 6416 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2157
timestamp 1018054153
transform 1 0 6432 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2159
timestamp 1018054153
transform 1 0 6448 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2161
timestamp 1018054153
transform 1 0 6464 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2163
timestamp 1018054153
transform 1 0 6480 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2165
timestamp 1018054153
transform 1 0 6496 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2167
timestamp 1018054153
transform 1 0 6512 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2169
timestamp 1018054153
transform 1 0 6528 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2171
timestamp 1018054153
transform 1 0 6544 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2173
timestamp 1018054153
transform 1 0 6560 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2175
timestamp 1018054153
transform 1 0 6576 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2177
timestamp 1018054153
transform 1 0 6592 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2179
timestamp 1018054153
transform 1 0 6608 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2181
timestamp 1018054153
transform 1 0 6624 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2183
timestamp 1018054153
transform 1 0 6640 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2185
timestamp 1018054153
transform 1 0 6656 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2187
timestamp 1018054153
transform 1 0 6672 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2189
timestamp 1018054153
transform 1 0 6688 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2191
timestamp 1018054153
transform 1 0 6704 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2193
timestamp 1018054153
transform 1 0 6720 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2195
timestamp 1018054153
transform 1 0 6736 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2197
timestamp 1018054153
transform 1 0 6752 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2199
timestamp 1018054153
transform 1 0 6768 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2201
timestamp 1018054153
transform 1 0 6784 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2203
timestamp 1018054153
transform 1 0 6800 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2205
timestamp 1018054153
transform 1 0 6816 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2207
timestamp 1018054153
transform 1 0 6832 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2209
timestamp 1018054153
transform 1 0 6848 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2211
timestamp 1018054153
transform 1 0 6864 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2213
timestamp 1018054153
transform 1 0 6880 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2215
timestamp 1018054153
transform 1 0 6896 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2217
timestamp 1018054153
transform 1 0 6912 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2219
timestamp 1018054153
transform 1 0 6928 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2221
timestamp 1018054153
transform 1 0 6944 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2223
timestamp 1018054153
transform 1 0 6960 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2225
timestamp 1018054153
transform 1 0 6976 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2227
timestamp 1018054153
transform 1 0 6992 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2229
timestamp 1018054153
transform 1 0 7008 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2231
timestamp 1018054153
transform 1 0 7024 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2233
timestamp 1018054153
transform 1 0 7040 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2235
timestamp 1018054153
transform 1 0 7056 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2237
timestamp 1018054153
transform 1 0 7072 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2239
timestamp 1018054153
transform 1 0 7088 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2241
timestamp 1018054153
transform 1 0 7104 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2243
timestamp 1018054153
transform 1 0 7120 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2245
timestamp 1018054153
transform 1 0 7136 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2247
timestamp 1018054153
transform 1 0 7152 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2249
timestamp 1018054153
transform 1 0 7168 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2251
timestamp 1018054153
transform 1 0 7184 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2253
timestamp 1018054153
transform 1 0 7200 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2255
timestamp 1018054153
transform 1 0 7216 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2257
timestamp 1018054153
transform 1 0 7232 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2259
timestamp 1018054153
transform 1 0 7248 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2261
timestamp 1018054153
transform 1 0 7264 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2263
timestamp 1018054153
transform 1 0 7280 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2265
timestamp 1018054153
transform 1 0 7296 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2267
timestamp 1018054153
transform 1 0 7312 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2269
timestamp 1018054153
transform 1 0 7328 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2271
timestamp 1018054153
transform 1 0 7344 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2273
timestamp 1018054153
transform 1 0 7360 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2275
timestamp 1018054153
transform 1 0 7376 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2277
timestamp 1018054153
transform 1 0 7392 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2279
timestamp 1018054153
transform 1 0 7408 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2281
timestamp 1018054153
transform 1 0 7424 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2283
timestamp 1018054153
transform 1 0 7440 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2285
timestamp 1018054153
transform 1 0 7456 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2287
timestamp 1018054153
transform 1 0 7472 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2289
timestamp 1018054153
transform 1 0 7488 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2291
timestamp 1018054153
transform 1 0 7504 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2293
timestamp 1018054153
transform 1 0 7520 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2295
timestamp 1018054153
transform 1 0 7536 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2297
timestamp 1018054153
transform 1 0 7552 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2299
timestamp 1018054153
transform 1 0 7568 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2301
timestamp 1018054153
transform 1 0 7584 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2303
timestamp 1018054153
transform 1 0 7600 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2305
timestamp 1018054153
transform 1 0 7616 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2307
timestamp 1018054153
transform 1 0 7632 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2309
timestamp 1018054153
transform 1 0 7648 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2311
timestamp 1018054153
transform 1 0 7664 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2313
timestamp 1018054153
transform 1 0 7680 0 -1 6480
box -16 -6 32 210
use FILL  FILL_2315
timestamp 1018054153
transform 1 0 7696 0 -1 6480
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_11
timestamp 1542725905
transform 1 0 7788 0 1 6280
box -48 -6 48 6
use FILL  FILL_2317
timestamp 1018054153
transform 1 0 7712 0 -1 6480
box -16 -6 32 210
use M2_M1  M2_M1_63
timestamp 1542725905
transform 1 0 3448 0 1 6170
box -4 -4 4 4
use M2_M1  M2_M1_70
timestamp 1542725905
transform 1 0 3432 0 1 6150
box -4 -4 4 4
use M2_M1  M2_M1_62
timestamp 1542725905
transform 1 0 3528 0 1 6190
box -4 -4 4 4
use M2_M1  M2_M1_71
timestamp 1542725905
transform 1 0 3816 0 1 6150
box -4 -4 4 4
use M3_M2  M3_M2_24
timestamp 1542725905
transform 1 0 3800 0 1 6130
box -6 -6 6 6
use M3_M2  M3_M2_21
timestamp 1542725905
transform 1 0 3832 0 1 6150
box -6 -6 6 6
use M2_M1  M2_M1_72
timestamp 1542725905
transform 1 0 3848 0 1 6150
box -4 -4 4 4
use M2_M1  M2_M1_78
timestamp 1542725905
transform 1 0 4056 0 1 6130
box -4 -4 4 4
use M2_M1  M2_M1_64
timestamp 1542725905
transform 1 0 4184 0 1 6170
box -4 -4 4 4
use M3_M2  M3_M2_25
timestamp 1542725905
transform 1 0 4344 0 1 6110
box -6 -6 6 6
use M2_M1  M2_M1_65
timestamp 1542725905
transform 1 0 4584 0 1 6170
box -4 -4 4 4
use M2_M1  M2_M1_73
timestamp 1542725905
transform 1 0 4712 0 1 6150
box -4 -4 4 4
use M3_M2  M3_M2_15
timestamp 1542725905
transform 1 0 4808 0 1 6210
box -6 -6 6 6
use M3_M2  M3_M2_16
timestamp 1542725905
transform 1 0 4920 0 1 6210
box -6 -6 6 6
use M2_M1  M2_M1_66
timestamp 1542725905
transform 1 0 4760 0 1 6170
box -4 -4 4 4
use M3_M2  M3_M2_17
timestamp 1542725905
transform 1 0 4808 0 1 6170
box -6 -6 6 6
use M2_M1  M2_M1_79
timestamp 1542725905
transform 1 0 4936 0 1 6130
box -4 -4 4 4
use M3_M2  M3_M2_26
timestamp 1542725905
transform 1 0 4744 0 1 6110
box -6 -6 6 6
use M3_M2  M3_M2_27
timestamp 1542725905
transform 1 0 4936 0 1 6110
box -6 -6 6 6
use M2_M1  M2_M1_67
timestamp 1542725905
transform 1 0 5176 0 1 6170
box -4 -4 4 4
use M2_M1  M2_M1_68
timestamp 1542725905
transform 1 0 5192 0 1 6170
box -4 -4 4 4
use M3_M2  M3_M2_18
timestamp 1542725905
transform 1 0 5256 0 1 6170
box -6 -6 6 6
use M3_M2  M3_M2_22
timestamp 1542725905
transform 1 0 5192 0 1 6150
box -6 -6 6 6
use M2_M1  M2_M1_80
timestamp 1542725905
transform 1 0 5368 0 1 6130
box -4 -4 4 4
use M3_M2  M3_M2_13
timestamp 1542725905
transform 1 0 5496 0 1 6250
box -6 -6 6 6
use M3_M2  M3_M2_28
timestamp 1542725905
transform 1 0 5480 0 1 6110
box -6 -6 6 6
use M2_M1  M2_M1_69
timestamp 1542725905
transform 1 0 5592 0 1 6170
box -4 -4 4 4
use M2_M1  M2_M1_74
timestamp 1542725905
transform 1 0 5608 0 1 6150
box -4 -4 4 4
use M3_M2  M3_M2_19
timestamp 1542725905
transform 1 0 5640 0 1 6170
box -6 -6 6 6
use M2_M1  M2_M1_75
timestamp 1542725905
transform 1 0 5640 0 1 6150
box -4 -4 4 4
use M2_M1  M2_M1_81
timestamp 1542725905
transform 1 0 5672 0 1 6130
box -4 -4 4 4
use M3_M2  M3_M2_20
timestamp 1542725905
transform 1 0 5768 0 1 6170
box -6 -6 6 6
use M2_M1  M2_M1_76
timestamp 1542725905
transform 1 0 5880 0 1 6150
box -4 -4 4 4
use M2_M1  M2_M1_82
timestamp 1542725905
transform 1 0 5944 0 1 6130
box -4 -4 4 4
use M3_M2  M3_M2_14
timestamp 1542725905
transform 1 0 5976 0 1 6250
box -6 -6 6 6
use M2_M1  M2_M1_83
timestamp 1542725905
transform 1 0 5976 0 1 6130
box -4 -4 4 4
use M2_M1  M2_M1_77
timestamp 1542725905
transform 1 0 6008 0 1 6150
box -4 -4 4 4
use PADNC  PADNC_6
timestamp 1084294400
transform 0 1 8000 -1 0 6800
box -6 -6 606 2000
use mult_pad_VIA1  mult_pad_VIA1_12
timestamp 1542725905
transform 1 0 2092 0 1 6080
box -48 -6 48 6
use FILL  FILL_2318
timestamp 1018054153
transform 1 0 2272 0 1 6080
box -16 -6 32 210
use FILL  FILL_2320
timestamp 1018054153
transform 1 0 2288 0 1 6080
box -16 -6 32 210
use FILL  FILL_2322
timestamp 1018054153
transform 1 0 2304 0 1 6080
box -16 -6 32 210
use FILL  FILL_2324
timestamp 1018054153
transform 1 0 2320 0 1 6080
box -16 -6 32 210
use FILL  FILL_2326
timestamp 1018054153
transform 1 0 2336 0 1 6080
box -16 -6 32 210
use FILL  FILL_2328
timestamp 1018054153
transform 1 0 2352 0 1 6080
box -16 -6 32 210
use FILL  FILL_2330
timestamp 1018054153
transform 1 0 2368 0 1 6080
box -16 -6 32 210
use FILL  FILL_2332
timestamp 1018054153
transform 1 0 2384 0 1 6080
box -16 -6 32 210
use FILL  FILL_2334
timestamp 1018054153
transform 1 0 2400 0 1 6080
box -16 -6 32 210
use FILL  FILL_2336
timestamp 1018054153
transform 1 0 2416 0 1 6080
box -16 -6 32 210
use FILL  FILL_2338
timestamp 1018054153
transform 1 0 2432 0 1 6080
box -16 -6 32 210
use FILL  FILL_2340
timestamp 1018054153
transform 1 0 2448 0 1 6080
box -16 -6 32 210
use FILL  FILL_2342
timestamp 1018054153
transform 1 0 2464 0 1 6080
box -16 -6 32 210
use FILL  FILL_2344
timestamp 1018054153
transform 1 0 2480 0 1 6080
box -16 -6 32 210
use FILL  FILL_2346
timestamp 1018054153
transform 1 0 2496 0 1 6080
box -16 -6 32 210
use FILL  FILL_2348
timestamp 1018054153
transform 1 0 2512 0 1 6080
box -16 -6 32 210
use FILL  FILL_2350
timestamp 1018054153
transform 1 0 2528 0 1 6080
box -16 -6 32 210
use FILL  FILL_2352
timestamp 1018054153
transform 1 0 2544 0 1 6080
box -16 -6 32 210
use FILL  FILL_2354
timestamp 1018054153
transform 1 0 2560 0 1 6080
box -16 -6 32 210
use FILL  FILL_2356
timestamp 1018054153
transform 1 0 2576 0 1 6080
box -16 -6 32 210
use FILL  FILL_2358
timestamp 1018054153
transform 1 0 2592 0 1 6080
box -16 -6 32 210
use FILL  FILL_2360
timestamp 1018054153
transform 1 0 2608 0 1 6080
box -16 -6 32 210
use FILL  FILL_2362
timestamp 1018054153
transform 1 0 2624 0 1 6080
box -16 -6 32 210
use FILL  FILL_2364
timestamp 1018054153
transform 1 0 2640 0 1 6080
box -16 -6 32 210
use FILL  FILL_2366
timestamp 1018054153
transform 1 0 2656 0 1 6080
box -16 -6 32 210
use FILL  FILL_2368
timestamp 1018054153
transform 1 0 2672 0 1 6080
box -16 -6 32 210
use FILL  FILL_2370
timestamp 1018054153
transform 1 0 2688 0 1 6080
box -16 -6 32 210
use FILL  FILL_2372
timestamp 1018054153
transform 1 0 2704 0 1 6080
box -16 -6 32 210
use FILL  FILL_2374
timestamp 1018054153
transform 1 0 2720 0 1 6080
box -16 -6 32 210
use FILL  FILL_2376
timestamp 1018054153
transform 1 0 2736 0 1 6080
box -16 -6 32 210
use FILL  FILL_2378
timestamp 1018054153
transform 1 0 2752 0 1 6080
box -16 -6 32 210
use FILL  FILL_2380
timestamp 1018054153
transform 1 0 2768 0 1 6080
box -16 -6 32 210
use FILL  FILL_2382
timestamp 1018054153
transform 1 0 2784 0 1 6080
box -16 -6 32 210
use FILL  FILL_2384
timestamp 1018054153
transform 1 0 2800 0 1 6080
box -16 -6 32 210
use FILL  FILL_2386
timestamp 1018054153
transform 1 0 2816 0 1 6080
box -16 -6 32 210
use FILL  FILL_2388
timestamp 1018054153
transform 1 0 2832 0 1 6080
box -16 -6 32 210
use FILL  FILL_2390
timestamp 1018054153
transform 1 0 2848 0 1 6080
box -16 -6 32 210
use FILL  FILL_2392
timestamp 1018054153
transform 1 0 2864 0 1 6080
box -16 -6 32 210
use FILL  FILL_2394
timestamp 1018054153
transform 1 0 2880 0 1 6080
box -16 -6 32 210
use FILL  FILL_2396
timestamp 1018054153
transform 1 0 2896 0 1 6080
box -16 -6 32 210
use FILL  FILL_2398
timestamp 1018054153
transform 1 0 2912 0 1 6080
box -16 -6 32 210
use FILL  FILL_2400
timestamp 1018054153
transform 1 0 2928 0 1 6080
box -16 -6 32 210
use FILL  FILL_2402
timestamp 1018054153
transform 1 0 2944 0 1 6080
box -16 -6 32 210
use FILL  FILL_2404
timestamp 1018054153
transform 1 0 2960 0 1 6080
box -16 -6 32 210
use FILL  FILL_2406
timestamp 1018054153
transform 1 0 2976 0 1 6080
box -16 -6 32 210
use FILL  FILL_2408
timestamp 1018054153
transform 1 0 2992 0 1 6080
box -16 -6 32 210
use FILL  FILL_2410
timestamp 1018054153
transform 1 0 3008 0 1 6080
box -16 -6 32 210
use FILL  FILL_2412
timestamp 1018054153
transform 1 0 3024 0 1 6080
box -16 -6 32 210
use FILL  FILL_2414
timestamp 1018054153
transform 1 0 3040 0 1 6080
box -16 -6 32 210
use FILL  FILL_2416
timestamp 1018054153
transform 1 0 3056 0 1 6080
box -16 -6 32 210
use FILL  FILL_2418
timestamp 1018054153
transform 1 0 3072 0 1 6080
box -16 -6 32 210
use FILL  FILL_2420
timestamp 1018054153
transform 1 0 3088 0 1 6080
box -16 -6 32 210
use FILL  FILL_2422
timestamp 1018054153
transform 1 0 3104 0 1 6080
box -16 -6 32 210
use FILL  FILL_2424
timestamp 1018054153
transform 1 0 3120 0 1 6080
box -16 -6 32 210
use FILL  FILL_2426
timestamp 1018054153
transform 1 0 3136 0 1 6080
box -16 -6 32 210
use FILL  FILL_2428
timestamp 1018054153
transform 1 0 3152 0 1 6080
box -16 -6 32 210
use FILL  FILL_2430
timestamp 1018054153
transform 1 0 3168 0 1 6080
box -16 -6 32 210
use FILL  FILL_2432
timestamp 1018054153
transform 1 0 3184 0 1 6080
box -16 -6 32 210
use FILL  FILL_2434
timestamp 1018054153
transform 1 0 3200 0 1 6080
box -16 -6 32 210
use FILL  FILL_2436
timestamp 1018054153
transform 1 0 3216 0 1 6080
box -16 -6 32 210
use FILL  FILL_2438
timestamp 1018054153
transform 1 0 3232 0 1 6080
box -16 -6 32 210
use FILL  FILL_2440
timestamp 1018054153
transform 1 0 3248 0 1 6080
box -16 -6 32 210
use FILL  FILL_2442
timestamp 1018054153
transform 1 0 3264 0 1 6080
box -16 -6 32 210
use FILL  FILL_2444
timestamp 1018054153
transform 1 0 3280 0 1 6080
box -16 -6 32 210
use FILL  FILL_2446
timestamp 1018054153
transform 1 0 3296 0 1 6080
box -16 -6 32 210
use FILL  FILL_2448
timestamp 1018054153
transform 1 0 3312 0 1 6080
box -16 -6 32 210
use FILL  FILL_2450
timestamp 1018054153
transform 1 0 3328 0 1 6080
box -16 -6 32 210
use FILL  FILL_2452
timestamp 1018054153
transform 1 0 3344 0 1 6080
box -16 -6 32 210
use FILL  FILL_2454
timestamp 1018054153
transform 1 0 3360 0 1 6080
box -16 -6 32 210
use FILL  FILL_2456
timestamp 1018054153
transform 1 0 3376 0 1 6080
box -16 -6 32 210
use FILL  FILL_2458
timestamp 1018054153
transform 1 0 3392 0 1 6080
box -16 -6 32 210
use FILL  FILL_2460
timestamp 1018054153
transform 1 0 3408 0 1 6080
box -16 -6 32 210
use OAI21X1  OAI21X1_7
timestamp 1053722159
transform 1 0 3424 0 1 6080
box -16 -6 68 210
use FILL  FILL_2462
timestamp 1018054153
transform 1 0 3488 0 1 6080
box -16 -6 32 210
use FILL  FILL_2468
timestamp 1018054153
transform 1 0 3504 0 1 6080
box -16 -6 32 210
use FILL  FILL_2470
timestamp 1018054153
transform 1 0 3520 0 1 6080
box -16 -6 32 210
use FILL  FILL_2472
timestamp 1018054153
transform 1 0 3536 0 1 6080
box -16 -6 32 210
use FILL  FILL_2474
timestamp 1018054153
transform 1 0 3552 0 1 6080
box -16 -6 32 210
use FILL  FILL_2476
timestamp 1018054153
transform 1 0 3568 0 1 6080
box -16 -6 32 210
use FILL  FILL_2478
timestamp 1018054153
transform 1 0 3584 0 1 6080
box -16 -6 32 210
use FILL  FILL_2480
timestamp 1018054153
transform 1 0 3600 0 1 6080
box -16 -6 32 210
use FILL  FILL_2482
timestamp 1018054153
transform 1 0 3616 0 1 6080
box -16 -6 32 210
use FILL  FILL_2484
timestamp 1018054153
transform 1 0 3632 0 1 6080
box -16 -6 32 210
use FILL  FILL_2486
timestamp 1018054153
transform 1 0 3648 0 1 6080
box -16 -6 32 210
use FILL  FILL_2488
timestamp 1018054153
transform 1 0 3664 0 1 6080
box -16 -6 32 210
use FILL  FILL_2490
timestamp 1018054153
transform 1 0 3680 0 1 6080
box -16 -6 32 210
use FILL  FILL_2492
timestamp 1018054153
transform 1 0 3696 0 1 6080
box -16 -6 32 210
use FILL  FILL_2494
timestamp 1018054153
transform 1 0 3712 0 1 6080
box -16 -6 32 210
use FILL  FILL_2496
timestamp 1018054153
transform 1 0 3728 0 1 6080
box -16 -6 32 210
use FILL  FILL_2498
timestamp 1018054153
transform 1 0 3744 0 1 6080
box -16 -6 32 210
use FILL  FILL_2500
timestamp 1018054153
transform 1 0 3760 0 1 6080
box -16 -6 32 210
use FILL  FILL_2502
timestamp 1018054153
transform 1 0 3776 0 1 6080
box -16 -6 32 210
use FILL  FILL_2504
timestamp 1018054153
transform 1 0 3792 0 1 6080
box -16 -6 32 210
use FILL  FILL_2506
timestamp 1018054153
transform 1 0 3808 0 1 6080
box -16 -6 32 210
use FILL  FILL_2508
timestamp 1018054153
transform 1 0 3824 0 1 6080
box -16 -6 32 210
use FILL  FILL_2510
timestamp 1018054153
transform 1 0 3840 0 1 6080
box -16 -6 32 210
use FILL  FILL_2512
timestamp 1018054153
transform 1 0 3856 0 1 6080
box -16 -6 32 210
use FILL  FILL_2514
timestamp 1018054153
transform 1 0 3872 0 1 6080
box -16 -6 32 210
use FILL  FILL_2516
timestamp 1018054153
transform 1 0 3888 0 1 6080
box -16 -6 32 210
use FILL  FILL_2518
timestamp 1018054153
transform 1 0 3904 0 1 6080
box -16 -6 32 210
use FILL  FILL_2520
timestamp 1018054153
transform 1 0 3920 0 1 6080
box -16 -6 32 210
use FILL  FILL_2522
timestamp 1018054153
transform 1 0 3936 0 1 6080
box -16 -6 32 210
use FILL  FILL_2524
timestamp 1018054153
transform 1 0 3952 0 1 6080
box -16 -6 32 210
use FILL  FILL_2526
timestamp 1018054153
transform 1 0 3968 0 1 6080
box -16 -6 32 210
use FILL  FILL_2527
timestamp 1018054153
transform 1 0 3984 0 1 6080
box -16 -6 32 210
use FILL  FILL_2528
timestamp 1018054153
transform 1 0 4000 0 1 6080
box -16 -6 32 210
use FILL  FILL_2529
timestamp 1018054153
transform 1 0 4016 0 1 6080
box -16 -6 32 210
use FILL  FILL_2530
timestamp 1018054153
transform 1 0 4032 0 1 6080
box -16 -6 32 210
use FILL  FILL_2531
timestamp 1018054153
transform 1 0 4048 0 1 6080
box -16 -6 32 210
use FILL  FILL_2534
timestamp 1018054153
transform 1 0 4064 0 1 6080
box -16 -6 32 210
use FILL  FILL_2536
timestamp 1018054153
transform 1 0 4080 0 1 6080
box -16 -6 32 210
use FILL  FILL_2538
timestamp 1018054153
transform 1 0 4096 0 1 6080
box -16 -6 32 210
use FILL  FILL_2540
timestamp 1018054153
transform 1 0 4112 0 1 6080
box -16 -6 32 210
use NOR2X1  NOR2X1_2
timestamp 1053022145
transform 1 0 4128 0 1 6080
box -16 -6 64 210
use FILL  FILL_2542
timestamp 1018054153
transform 1 0 4176 0 1 6080
box -16 -6 32 210
use FILL  FILL_2547
timestamp 1018054153
transform 1 0 4192 0 1 6080
box -16 -6 32 210
use FILL  FILL_2549
timestamp 1018054153
transform 1 0 4208 0 1 6080
box -16 -6 32 210
use FILL  FILL_2551
timestamp 1018054153
transform 1 0 4224 0 1 6080
box -16 -6 32 210
use FILL  FILL_2553
timestamp 1018054153
transform 1 0 4240 0 1 6080
box -16 -6 32 210
use FILL  FILL_2555
timestamp 1018054153
transform 1 0 4256 0 1 6080
box -16 -6 32 210
use FILL  FILL_2557
timestamp 1018054153
transform 1 0 4272 0 1 6080
box -16 -6 32 210
use FILL  FILL_2559
timestamp 1018054153
transform 1 0 4288 0 1 6080
box -16 -6 32 210
use FILL  FILL_2561
timestamp 1018054153
transform 1 0 4304 0 1 6080
box -16 -6 32 210
use FILL  FILL_2563
timestamp 1018054153
transform 1 0 4320 0 1 6080
box -16 -6 32 210
use FILL  FILL_2565
timestamp 1018054153
transform 1 0 4336 0 1 6080
box -16 -6 32 210
use FILL  FILL_2567
timestamp 1018054153
transform 1 0 4352 0 1 6080
box -16 -6 32 210
use FILL  FILL_2569
timestamp 1018054153
transform 1 0 4368 0 1 6080
box -16 -6 32 210
use FILL  FILL_2571
timestamp 1018054153
transform 1 0 4384 0 1 6080
box -16 -6 32 210
use FILL  FILL_2573
timestamp 1018054153
transform 1 0 4400 0 1 6080
box -16 -6 32 210
use FILL  FILL_2575
timestamp 1018054153
transform 1 0 4416 0 1 6080
box -16 -6 32 210
use FILL  FILL_2577
timestamp 1018054153
transform 1 0 4432 0 1 6080
box -16 -6 32 210
use FILL  FILL_2579
timestamp 1018054153
transform 1 0 4448 0 1 6080
box -16 -6 32 210
use FILL  FILL_2581
timestamp 1018054153
transform 1 0 4464 0 1 6080
box -16 -6 32 210
use FILL  FILL_2583
timestamp 1018054153
transform 1 0 4480 0 1 6080
box -16 -6 32 210
use FILL  FILL_2585
timestamp 1018054153
transform 1 0 4496 0 1 6080
box -16 -6 32 210
use FILL  FILL_2586
timestamp 1018054153
transform 1 0 4512 0 1 6080
box -16 -6 32 210
use FILL  FILL_2587
timestamp 1018054153
transform 1 0 4528 0 1 6080
box -16 -6 32 210
use FILL  FILL_2588
timestamp 1018054153
transform 1 0 4544 0 1 6080
box -16 -6 32 210
use FILL  FILL_2590
timestamp 1018054153
transform 1 0 4560 0 1 6080
box -16 -6 32 210
use FILL  FILL_2592
timestamp 1018054153
transform 1 0 4576 0 1 6080
box -16 -6 32 210
use FILL  FILL_2594
timestamp 1018054153
transform 1 0 4592 0 1 6080
box -16 -6 32 210
use FILL  FILL_2596
timestamp 1018054153
transform 1 0 4608 0 1 6080
box -16 -6 32 210
use FILL  FILL_2598
timestamp 1018054153
transform 1 0 4624 0 1 6080
box -16 -6 32 210
use FILL  FILL_2600
timestamp 1018054153
transform 1 0 4640 0 1 6080
box -16 -6 32 210
use FILL  FILL_2602
timestamp 1018054153
transform 1 0 4656 0 1 6080
box -16 -6 32 210
use FILL  FILL_2604
timestamp 1018054153
transform 1 0 4672 0 1 6080
box -16 -6 32 210
use FILL  FILL_2606
timestamp 1018054153
transform 1 0 4688 0 1 6080
box -16 -6 32 210
use FILL  FILL_2608
timestamp 1018054153
transform 1 0 4704 0 1 6080
box -16 -6 32 210
use FAX1  FAX1_0
timestamp 1053025068
transform 1 0 4720 0 1 6080
box -10 -6 252 210
use FILL  FILL_2610
timestamp 1018054153
transform 1 0 4960 0 1 6080
box -16 -6 32 210
use FILL  FILL_2624
timestamp 1018054153
transform 1 0 4976 0 1 6080
box -16 -6 32 210
use FILL  FILL_2626
timestamp 1018054153
transform 1 0 4992 0 1 6080
box -16 -6 32 210
use FILL  FILL_2628
timestamp 1018054153
transform 1 0 5008 0 1 6080
box -16 -6 32 210
use FILL  FILL_2630
timestamp 1018054153
transform 1 0 5024 0 1 6080
box -16 -6 32 210
use FILL  FILL_2632
timestamp 1018054153
transform 1 0 5040 0 1 6080
box -16 -6 32 210
use FILL  FILL_2634
timestamp 1018054153
transform 1 0 5056 0 1 6080
box -16 -6 32 210
use FILL  FILL_2636
timestamp 1018054153
transform 1 0 5072 0 1 6080
box -16 -6 32 210
use FILL  FILL_2638
timestamp 1018054153
transform 1 0 5088 0 1 6080
box -16 -6 32 210
use FILL  FILL_2640
timestamp 1018054153
transform 1 0 5104 0 1 6080
box -16 -6 32 210
use FILL  FILL_2642
timestamp 1018054153
transform 1 0 5120 0 1 6080
box -16 -6 32 210
use FILL  FILL_2644
timestamp 1018054153
transform 1 0 5136 0 1 6080
box -16 -6 32 210
use FAX1  FAX1_1
timestamp 1053025068
transform 1 0 5152 0 1 6080
box -10 -6 252 210
use FILL  FILL_2646
timestamp 1018054153
transform 1 0 5392 0 1 6080
box -16 -6 32 210
use FILL  FILL_2660
timestamp 1018054153
transform 1 0 5408 0 1 6080
box -16 -6 32 210
use FILL  FILL_2662
timestamp 1018054153
transform 1 0 5424 0 1 6080
box -16 -6 32 210
use FILL  FILL_2664
timestamp 1018054153
transform 1 0 5440 0 1 6080
box -16 -6 32 210
use FILL  FILL_2666
timestamp 1018054153
transform 1 0 5456 0 1 6080
box -16 -6 32 210
use FILL  FILL_2668
timestamp 1018054153
transform 1 0 5472 0 1 6080
box -16 -6 32 210
use FILL  FILL_2670
timestamp 1018054153
transform 1 0 5488 0 1 6080
box -16 -6 32 210
use FILL  FILL_2672
timestamp 1018054153
transform 1 0 5504 0 1 6080
box -16 -6 32 210
use FILL  FILL_2674
timestamp 1018054153
transform 1 0 5520 0 1 6080
box -16 -6 32 210
use FILL  FILL_2676
timestamp 1018054153
transform 1 0 5536 0 1 6080
box -16 -6 32 210
use FILL  FILL_2678
timestamp 1018054153
transform 1 0 5552 0 1 6080
box -16 -6 32 210
use FILL  FILL_2680
timestamp 1018054153
transform 1 0 5568 0 1 6080
box -16 -6 32 210
use FILL  FILL_2682
timestamp 1018054153
transform 1 0 5584 0 1 6080
box -16 -6 32 210
use FILL  FILL_2684
timestamp 1018054153
transform 1 0 5600 0 1 6080
box -16 -6 32 210
use AOI21X1  AOI21X1_0
timestamp 1090541997
transform 1 0 5616 0 1 6080
box -14 -6 78 210
use FILL  FILL_2686
timestamp 1018054153
transform 1 0 5680 0 1 6080
box -16 -6 32 210
use FILL  FILL_2687
timestamp 1018054153
transform 1 0 5696 0 1 6080
box -16 -6 32 210
use FILL  FILL_2688
timestamp 1018054153
transform 1 0 5712 0 1 6080
box -16 -6 32 210
use FILL  FILL_2689
timestamp 1018054153
transform 1 0 5728 0 1 6080
box -16 -6 32 210
use FILL  FILL_2690
timestamp 1018054153
transform 1 0 5744 0 1 6080
box -16 -6 32 210
use FILL  FILL_2691
timestamp 1018054153
transform 1 0 5760 0 1 6080
box -16 -6 32 210
use FILL  FILL_2692
timestamp 1018054153
transform 1 0 5776 0 1 6080
box -16 -6 32 210
use FILL  FILL_2697
timestamp 1018054153
transform 1 0 5792 0 1 6080
box -16 -6 32 210
use FILL  FILL_2699
timestamp 1018054153
transform 1 0 5808 0 1 6080
box -16 -6 32 210
use FILL  FILL_2701
timestamp 1018054153
transform 1 0 5824 0 1 6080
box -16 -6 32 210
use FILL  FILL_2703
timestamp 1018054153
transform 1 0 5840 0 1 6080
box -16 -6 32 210
use FILL  FILL_2705
timestamp 1018054153
transform 1 0 5856 0 1 6080
box -16 -6 32 210
use FILL  FILL_2707
timestamp 1018054153
transform 1 0 5872 0 1 6080
box -16 -6 32 210
use FILL  FILL_2709
timestamp 1018054153
transform 1 0 5888 0 1 6080
box -16 -6 32 210
use FILL  FILL_2711
timestamp 1018054153
transform 1 0 5904 0 1 6080
box -16 -6 32 210
use FILL  FILL_2713
timestamp 1018054153
transform 1 0 5920 0 1 6080
box -16 -6 32 210
use FILL  FILL_2715
timestamp 1018054153
transform 1 0 5936 0 1 6080
box -16 -6 32 210
use FILL  FILL_2717
timestamp 1018054153
transform 1 0 5952 0 1 6080
box -16 -6 32 210
use FILL  FILL_2718
timestamp 1018054153
transform 1 0 5968 0 1 6080
box -16 -6 32 210
use FILL  FILL_2719
timestamp 1018054153
transform 1 0 5984 0 1 6080
box -16 -6 32 210
use FILL  FILL_2720
timestamp 1018054153
transform 1 0 6000 0 1 6080
box -16 -6 32 210
use FILL  FILL_2721
timestamp 1018054153
transform 1 0 6016 0 1 6080
box -16 -6 32 210
use FILL  FILL_2723
timestamp 1018054153
transform 1 0 6032 0 1 6080
box -16 -6 32 210
use FILL  FILL_2725
timestamp 1018054153
transform 1 0 6048 0 1 6080
box -16 -6 32 210
use FILL  FILL_2727
timestamp 1018054153
transform 1 0 6064 0 1 6080
box -16 -6 32 210
use FILL  FILL_2729
timestamp 1018054153
transform 1 0 6080 0 1 6080
box -16 -6 32 210
use FILL  FILL_2731
timestamp 1018054153
transform 1 0 6096 0 1 6080
box -16 -6 32 210
use FILL  FILL_2733
timestamp 1018054153
transform 1 0 6112 0 1 6080
box -16 -6 32 210
use FILL  FILL_2735
timestamp 1018054153
transform 1 0 6128 0 1 6080
box -16 -6 32 210
use FILL  FILL_2737
timestamp 1018054153
transform 1 0 6144 0 1 6080
box -16 -6 32 210
use FILL  FILL_2739
timestamp 1018054153
transform 1 0 6160 0 1 6080
box -16 -6 32 210
use FILL  FILL_2741
timestamp 1018054153
transform 1 0 6176 0 1 6080
box -16 -6 32 210
use FILL  FILL_2743
timestamp 1018054153
transform 1 0 6192 0 1 6080
box -16 -6 32 210
use INVX1  INVX1_5
timestamp 1053022145
transform 1 0 6208 0 1 6080
box -18 -6 52 210
use FILL  FILL_2745
timestamp 1018054153
transform 1 0 6240 0 1 6080
box -16 -6 32 210
use FILL  FILL_2749
timestamp 1018054153
transform 1 0 6256 0 1 6080
box -16 -6 32 210
use FILL  FILL_2751
timestamp 1018054153
transform 1 0 6272 0 1 6080
box -16 -6 32 210
use FILL  FILL_2753
timestamp 1018054153
transform 1 0 6288 0 1 6080
box -16 -6 32 210
use FILL  FILL_2755
timestamp 1018054153
transform 1 0 6304 0 1 6080
box -16 -6 32 210
use FILL  FILL_2757
timestamp 1018054153
transform 1 0 6320 0 1 6080
box -16 -6 32 210
use FILL  FILL_2759
timestamp 1018054153
transform 1 0 6336 0 1 6080
box -16 -6 32 210
use FILL  FILL_2761
timestamp 1018054153
transform 1 0 6352 0 1 6080
box -16 -6 32 210
use FILL  FILL_2763
timestamp 1018054153
transform 1 0 6368 0 1 6080
box -16 -6 32 210
use FILL  FILL_2765
timestamp 1018054153
transform 1 0 6384 0 1 6080
box -16 -6 32 210
use FILL  FILL_2767
timestamp 1018054153
transform 1 0 6400 0 1 6080
box -16 -6 32 210
use FILL  FILL_2769
timestamp 1018054153
transform 1 0 6416 0 1 6080
box -16 -6 32 210
use FILL  FILL_2771
timestamp 1018054153
transform 1 0 6432 0 1 6080
box -16 -6 32 210
use FILL  FILL_2773
timestamp 1018054153
transform 1 0 6448 0 1 6080
box -16 -6 32 210
use FILL  FILL_2775
timestamp 1018054153
transform 1 0 6464 0 1 6080
box -16 -6 32 210
use FILL  FILL_2777
timestamp 1018054153
transform 1 0 6480 0 1 6080
box -16 -6 32 210
use FILL  FILL_2779
timestamp 1018054153
transform 1 0 6496 0 1 6080
box -16 -6 32 210
use FILL  FILL_2781
timestamp 1018054153
transform 1 0 6512 0 1 6080
box -16 -6 32 210
use FILL  FILL_2783
timestamp 1018054153
transform 1 0 6528 0 1 6080
box -16 -6 32 210
use FILL  FILL_2785
timestamp 1018054153
transform 1 0 6544 0 1 6080
box -16 -6 32 210
use FILL  FILL_2787
timestamp 1018054153
transform 1 0 6560 0 1 6080
box -16 -6 32 210
use FILL  FILL_2789
timestamp 1018054153
transform 1 0 6576 0 1 6080
box -16 -6 32 210
use FILL  FILL_2791
timestamp 1018054153
transform 1 0 6592 0 1 6080
box -16 -6 32 210
use FILL  FILL_2793
timestamp 1018054153
transform 1 0 6608 0 1 6080
box -16 -6 32 210
use FILL  FILL_2795
timestamp 1018054153
transform 1 0 6624 0 1 6080
box -16 -6 32 210
use FILL  FILL_2797
timestamp 1018054153
transform 1 0 6640 0 1 6080
box -16 -6 32 210
use FILL  FILL_2799
timestamp 1018054153
transform 1 0 6656 0 1 6080
box -16 -6 32 210
use FILL  FILL_2801
timestamp 1018054153
transform 1 0 6672 0 1 6080
box -16 -6 32 210
use FILL  FILL_2803
timestamp 1018054153
transform 1 0 6688 0 1 6080
box -16 -6 32 210
use FILL  FILL_2805
timestamp 1018054153
transform 1 0 6704 0 1 6080
box -16 -6 32 210
use FILL  FILL_2807
timestamp 1018054153
transform 1 0 6720 0 1 6080
box -16 -6 32 210
use FILL  FILL_2809
timestamp 1018054153
transform 1 0 6736 0 1 6080
box -16 -6 32 210
use FILL  FILL_2811
timestamp 1018054153
transform 1 0 6752 0 1 6080
box -16 -6 32 210
use FILL  FILL_2813
timestamp 1018054153
transform 1 0 6768 0 1 6080
box -16 -6 32 210
use FILL  FILL_2815
timestamp 1018054153
transform 1 0 6784 0 1 6080
box -16 -6 32 210
use FILL  FILL_2817
timestamp 1018054153
transform 1 0 6800 0 1 6080
box -16 -6 32 210
use FILL  FILL_2819
timestamp 1018054153
transform 1 0 6816 0 1 6080
box -16 -6 32 210
use FILL  FILL_2821
timestamp 1018054153
transform 1 0 6832 0 1 6080
box -16 -6 32 210
use FILL  FILL_2823
timestamp 1018054153
transform 1 0 6848 0 1 6080
box -16 -6 32 210
use FILL  FILL_2825
timestamp 1018054153
transform 1 0 6864 0 1 6080
box -16 -6 32 210
use FILL  FILL_2827
timestamp 1018054153
transform 1 0 6880 0 1 6080
box -16 -6 32 210
use FILL  FILL_2829
timestamp 1018054153
transform 1 0 6896 0 1 6080
box -16 -6 32 210
use FILL  FILL_2831
timestamp 1018054153
transform 1 0 6912 0 1 6080
box -16 -6 32 210
use FILL  FILL_2833
timestamp 1018054153
transform 1 0 6928 0 1 6080
box -16 -6 32 210
use FILL  FILL_2835
timestamp 1018054153
transform 1 0 6944 0 1 6080
box -16 -6 32 210
use FILL  FILL_2837
timestamp 1018054153
transform 1 0 6960 0 1 6080
box -16 -6 32 210
use FILL  FILL_2839
timestamp 1018054153
transform 1 0 6976 0 1 6080
box -16 -6 32 210
use FILL  FILL_2841
timestamp 1018054153
transform 1 0 6992 0 1 6080
box -16 -6 32 210
use FILL  FILL_2843
timestamp 1018054153
transform 1 0 7008 0 1 6080
box -16 -6 32 210
use FILL  FILL_2845
timestamp 1018054153
transform 1 0 7024 0 1 6080
box -16 -6 32 210
use FILL  FILL_2847
timestamp 1018054153
transform 1 0 7040 0 1 6080
box -16 -6 32 210
use FILL  FILL_2849
timestamp 1018054153
transform 1 0 7056 0 1 6080
box -16 -6 32 210
use FILL  FILL_2851
timestamp 1018054153
transform 1 0 7072 0 1 6080
box -16 -6 32 210
use FILL  FILL_2853
timestamp 1018054153
transform 1 0 7088 0 1 6080
box -16 -6 32 210
use FILL  FILL_2855
timestamp 1018054153
transform 1 0 7104 0 1 6080
box -16 -6 32 210
use FILL  FILL_2857
timestamp 1018054153
transform 1 0 7120 0 1 6080
box -16 -6 32 210
use FILL  FILL_2859
timestamp 1018054153
transform 1 0 7136 0 1 6080
box -16 -6 32 210
use FILL  FILL_2861
timestamp 1018054153
transform 1 0 7152 0 1 6080
box -16 -6 32 210
use FILL  FILL_2863
timestamp 1018054153
transform 1 0 7168 0 1 6080
box -16 -6 32 210
use FILL  FILL_2865
timestamp 1018054153
transform 1 0 7184 0 1 6080
box -16 -6 32 210
use FILL  FILL_2867
timestamp 1018054153
transform 1 0 7200 0 1 6080
box -16 -6 32 210
use FILL  FILL_2869
timestamp 1018054153
transform 1 0 7216 0 1 6080
box -16 -6 32 210
use FILL  FILL_2871
timestamp 1018054153
transform 1 0 7232 0 1 6080
box -16 -6 32 210
use FILL  FILL_2873
timestamp 1018054153
transform 1 0 7248 0 1 6080
box -16 -6 32 210
use FILL  FILL_2875
timestamp 1018054153
transform 1 0 7264 0 1 6080
box -16 -6 32 210
use FILL  FILL_2877
timestamp 1018054153
transform 1 0 7280 0 1 6080
box -16 -6 32 210
use FILL  FILL_2879
timestamp 1018054153
transform 1 0 7296 0 1 6080
box -16 -6 32 210
use FILL  FILL_2881
timestamp 1018054153
transform 1 0 7312 0 1 6080
box -16 -6 32 210
use FILL  FILL_2883
timestamp 1018054153
transform 1 0 7328 0 1 6080
box -16 -6 32 210
use FILL  FILL_2885
timestamp 1018054153
transform 1 0 7344 0 1 6080
box -16 -6 32 210
use FILL  FILL_2887
timestamp 1018054153
transform 1 0 7360 0 1 6080
box -16 -6 32 210
use FILL  FILL_2889
timestamp 1018054153
transform 1 0 7376 0 1 6080
box -16 -6 32 210
use FILL  FILL_2891
timestamp 1018054153
transform 1 0 7392 0 1 6080
box -16 -6 32 210
use FILL  FILL_2893
timestamp 1018054153
transform 1 0 7408 0 1 6080
box -16 -6 32 210
use FILL  FILL_2895
timestamp 1018054153
transform 1 0 7424 0 1 6080
box -16 -6 32 210
use FILL  FILL_2897
timestamp 1018054153
transform 1 0 7440 0 1 6080
box -16 -6 32 210
use FILL  FILL_2899
timestamp 1018054153
transform 1 0 7456 0 1 6080
box -16 -6 32 210
use FILL  FILL_2901
timestamp 1018054153
transform 1 0 7472 0 1 6080
box -16 -6 32 210
use FILL  FILL_2903
timestamp 1018054153
transform 1 0 7488 0 1 6080
box -16 -6 32 210
use FILL  FILL_2905
timestamp 1018054153
transform 1 0 7504 0 1 6080
box -16 -6 32 210
use FILL  FILL_2907
timestamp 1018054153
transform 1 0 7520 0 1 6080
box -16 -6 32 210
use FILL  FILL_2909
timestamp 1018054153
transform 1 0 7536 0 1 6080
box -16 -6 32 210
use FILL  FILL_2911
timestamp 1018054153
transform 1 0 7552 0 1 6080
box -16 -6 32 210
use FILL  FILL_2913
timestamp 1018054153
transform 1 0 7568 0 1 6080
box -16 -6 32 210
use FILL  FILL_2915
timestamp 1018054153
transform 1 0 7584 0 1 6080
box -16 -6 32 210
use FILL  FILL_2917
timestamp 1018054153
transform 1 0 7600 0 1 6080
box -16 -6 32 210
use FILL  FILL_2919
timestamp 1018054153
transform 1 0 7616 0 1 6080
box -16 -6 32 210
use FILL  FILL_2921
timestamp 1018054153
transform 1 0 7632 0 1 6080
box -16 -6 32 210
use FILL  FILL_2923
timestamp 1018054153
transform 1 0 7648 0 1 6080
box -16 -6 32 210
use FILL  FILL_2925
timestamp 1018054153
transform 1 0 7664 0 1 6080
box -16 -6 32 210
use FILL  FILL_2927
timestamp 1018054153
transform 1 0 7680 0 1 6080
box -16 -6 32 210
use FILL  FILL_2929
timestamp 1018054153
transform 1 0 7696 0 1 6080
box -16 -6 32 210
use FILL  FILL_2931
timestamp 1018054153
transform 1 0 7712 0 1 6080
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_13
timestamp 1542725905
transform 1 0 7908 0 1 6080
box -48 -6 48 6
use M2_M1  M2_M1_85
timestamp 1542725905
transform 1 0 3512 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_100
timestamp 1542725905
transform 1 0 3912 0 1 5970
box -4 -4 4 4
use M2_M1  M2_M1_86
timestamp 1542725905
transform 1 0 4056 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_93
timestamp 1542725905
transform 1 0 4184 0 1 5990
box -4 -4 4 4
use M2_M1  M2_M1_87
timestamp 1542725905
transform 1 0 4456 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_103
timestamp 1542725905
transform 1 0 4552 0 1 5950
box -4 -4 4 4
use M2_M1  M2_M1_88
timestamp 1542725905
transform 1 0 4712 0 1 6010
box -4 -4 4 4
use M3_M2  M3_M2_32
timestamp 1542725905
transform 1 0 4808 0 1 6010
box -6 -6 6 6
use M2_M1  M2_M1_94
timestamp 1542725905
transform 1 0 4888 0 1 5990
box -4 -4 4 4
use M3_M2  M3_M2_35
timestamp 1542725905
transform 1 0 4888 0 1 5970
box -6 -6 6 6
use M2_M1  M2_M1_84
timestamp 1542725905
transform 1 0 4920 0 1 6030
box -4 -4 4 4
use M2_M1  M2_M1_95
timestamp 1542725905
transform 1 0 4968 0 1 5990
box -4 -4 4 4
use M3_M2  M3_M2_36
timestamp 1542725905
transform 1 0 4968 0 1 5970
box -6 -6 6 6
use M3_M2  M3_M2_33
timestamp 1542725905
transform 1 0 5128 0 1 6010
box -6 -6 6 6
use M2_M1  M2_M1_89
timestamp 1542725905
transform 1 0 5176 0 1 6010
box -4 -4 4 4
use M3_M2  M3_M2_34
timestamp 1542725905
transform 1 0 5320 0 1 6010
box -6 -6 6 6
use M2_M1  M2_M1_96
timestamp 1542725905
transform 1 0 5320 0 1 5990
box -4 -4 4 4
use M2_M1  M2_M1_90
timestamp 1542725905
transform 1 0 5384 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_97
timestamp 1542725905
transform 1 0 5368 0 1 5990
box -4 -4 4 4
use M3_M2  M3_M2_29
timestamp 1542725905
transform 1 0 5432 0 1 6070
box -6 -6 6 6
use M3_M2  M3_M2_30
timestamp 1542725905
transform 1 0 5592 0 1 6030
box -6 -6 6 6
use M2_M1  M2_M1_91
timestamp 1542725905
transform 1 0 5592 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_92
timestamp 1542725905
transform 1 0 5768 0 1 6010
box -4 -4 4 4
use M2_M1  M2_M1_98
timestamp 1542725905
transform 1 0 5736 0 1 5990
box -4 -4 4 4
use M2_M1  M2_M1_101
timestamp 1542725905
transform 1 0 5944 0 1 5970
box -4 -4 4 4
use M3_M2  M3_M2_31
timestamp 1542725905
transform 1 0 5976 0 1 6030
box -6 -6 6 6
use M2_M1  M2_M1_99
timestamp 1542725905
transform 1 0 5976 0 1 5990
box -4 -4 4 4
use M2_M1  M2_M1_102
timestamp 1542725905
transform 1 0 6024 0 1 5970
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_14
timestamp 1542725905
transform 1 0 2212 0 1 5880
box -48 -6 48 6
use FILL  FILL_2319
timestamp 1018054153
transform 1 0 2272 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2321
timestamp 1018054153
transform 1 0 2288 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2323
timestamp 1018054153
transform 1 0 2304 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2325
timestamp 1018054153
transform 1 0 2320 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2327
timestamp 1018054153
transform 1 0 2336 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2329
timestamp 1018054153
transform 1 0 2352 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2331
timestamp 1018054153
transform 1 0 2368 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2333
timestamp 1018054153
transform 1 0 2384 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2335
timestamp 1018054153
transform 1 0 2400 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2337
timestamp 1018054153
transform 1 0 2416 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2339
timestamp 1018054153
transform 1 0 2432 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2341
timestamp 1018054153
transform 1 0 2448 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2343
timestamp 1018054153
transform 1 0 2464 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2345
timestamp 1018054153
transform 1 0 2480 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2347
timestamp 1018054153
transform 1 0 2496 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2349
timestamp 1018054153
transform 1 0 2512 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2351
timestamp 1018054153
transform 1 0 2528 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2353
timestamp 1018054153
transform 1 0 2544 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2355
timestamp 1018054153
transform 1 0 2560 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2357
timestamp 1018054153
transform 1 0 2576 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2359
timestamp 1018054153
transform 1 0 2592 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2361
timestamp 1018054153
transform 1 0 2608 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2363
timestamp 1018054153
transform 1 0 2624 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2365
timestamp 1018054153
transform 1 0 2640 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2367
timestamp 1018054153
transform 1 0 2656 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2369
timestamp 1018054153
transform 1 0 2672 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2371
timestamp 1018054153
transform 1 0 2688 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2373
timestamp 1018054153
transform 1 0 2704 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2375
timestamp 1018054153
transform 1 0 2720 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2377
timestamp 1018054153
transform 1 0 2736 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2379
timestamp 1018054153
transform 1 0 2752 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2381
timestamp 1018054153
transform 1 0 2768 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2383
timestamp 1018054153
transform 1 0 2784 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2385
timestamp 1018054153
transform 1 0 2800 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2387
timestamp 1018054153
transform 1 0 2816 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2389
timestamp 1018054153
transform 1 0 2832 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2391
timestamp 1018054153
transform 1 0 2848 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2393
timestamp 1018054153
transform 1 0 2864 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2395
timestamp 1018054153
transform 1 0 2880 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2397
timestamp 1018054153
transform 1 0 2896 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2399
timestamp 1018054153
transform 1 0 2912 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2401
timestamp 1018054153
transform 1 0 2928 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2403
timestamp 1018054153
transform 1 0 2944 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2405
timestamp 1018054153
transform 1 0 2960 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2407
timestamp 1018054153
transform 1 0 2976 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2409
timestamp 1018054153
transform 1 0 2992 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2411
timestamp 1018054153
transform 1 0 3008 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2413
timestamp 1018054153
transform 1 0 3024 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2415
timestamp 1018054153
transform 1 0 3040 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2417
timestamp 1018054153
transform 1 0 3056 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2419
timestamp 1018054153
transform 1 0 3072 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2421
timestamp 1018054153
transform 1 0 3088 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2423
timestamp 1018054153
transform 1 0 3104 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2425
timestamp 1018054153
transform 1 0 3120 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2427
timestamp 1018054153
transform 1 0 3136 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2429
timestamp 1018054153
transform 1 0 3152 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2431
timestamp 1018054153
transform 1 0 3168 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2433
timestamp 1018054153
transform 1 0 3184 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2435
timestamp 1018054153
transform 1 0 3200 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2437
timestamp 1018054153
transform 1 0 3216 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2439
timestamp 1018054153
transform 1 0 3232 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2441
timestamp 1018054153
transform 1 0 3248 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2443
timestamp 1018054153
transform 1 0 3264 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2445
timestamp 1018054153
transform 1 0 3280 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2447
timestamp 1018054153
transform 1 0 3296 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2449
timestamp 1018054153
transform 1 0 3312 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2451
timestamp 1018054153
transform 1 0 3328 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2453
timestamp 1018054153
transform 1 0 3344 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2455
timestamp 1018054153
transform 1 0 3360 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2457
timestamp 1018054153
transform 1 0 3376 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2459
timestamp 1018054153
transform 1 0 3392 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2461
timestamp 1018054153
transform 1 0 3408 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2463
timestamp 1018054153
transform 1 0 3424 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2464
timestamp 1018054153
transform 1 0 3440 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2465
timestamp 1018054153
transform 1 0 3456 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2466
timestamp 1018054153
transform 1 0 3472 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2467
timestamp 1018054153
transform 1 0 3488 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2469
timestamp 1018054153
transform 1 0 3504 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2471
timestamp 1018054153
transform 1 0 3520 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2473
timestamp 1018054153
transform 1 0 3536 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2475
timestamp 1018054153
transform 1 0 3552 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2477
timestamp 1018054153
transform 1 0 3568 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2479
timestamp 1018054153
transform 1 0 3584 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2481
timestamp 1018054153
transform 1 0 3600 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2483
timestamp 1018054153
transform 1 0 3616 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2485
timestamp 1018054153
transform 1 0 3632 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2487
timestamp 1018054153
transform 1 0 3648 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2489
timestamp 1018054153
transform 1 0 3664 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2491
timestamp 1018054153
transform 1 0 3680 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2493
timestamp 1018054153
transform 1 0 3696 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2495
timestamp 1018054153
transform 1 0 3712 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2497
timestamp 1018054153
transform 1 0 3728 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2499
timestamp 1018054153
transform 1 0 3744 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2501
timestamp 1018054153
transform 1 0 3760 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2503
timestamp 1018054153
transform 1 0 3776 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2505
timestamp 1018054153
transform 1 0 3792 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2507
timestamp 1018054153
transform 1 0 3808 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2509
timestamp 1018054153
transform 1 0 3824 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2511
timestamp 1018054153
transform 1 0 3840 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2513
timestamp 1018054153
transform 1 0 3856 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2515
timestamp 1018054153
transform 1 0 3872 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2517
timestamp 1018054153
transform 1 0 3888 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2519
timestamp 1018054153
transform 1 0 3904 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2521
timestamp 1018054153
transform 1 0 3920 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2523
timestamp 1018054153
transform 1 0 3936 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2525
timestamp 1018054153
transform 1 0 3952 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2532
timestamp 1018054153
transform 1 0 3968 0 -1 6080
box -16 -6 32 210
use OAI21X1  OAI21X1_8
timestamp 1053722159
transform -1 0 4048 0 -1 6080
box -16 -6 68 210
use FILL  FILL_2533
timestamp 1018054153
transform 1 0 4048 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2535
timestamp 1018054153
transform 1 0 4064 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2537
timestamp 1018054153
transform 1 0 4080 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2539
timestamp 1018054153
transform 1 0 4096 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2541
timestamp 1018054153
transform 1 0 4112 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2543
timestamp 1018054153
transform 1 0 4128 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2544
timestamp 1018054153
transform 1 0 4144 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2545
timestamp 1018054153
transform 1 0 4160 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2546
timestamp 1018054153
transform 1 0 4176 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2548
timestamp 1018054153
transform 1 0 4192 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2550
timestamp 1018054153
transform 1 0 4208 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2552
timestamp 1018054153
transform 1 0 4224 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2554
timestamp 1018054153
transform 1 0 4240 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2556
timestamp 1018054153
transform 1 0 4256 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2558
timestamp 1018054153
transform 1 0 4272 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2560
timestamp 1018054153
transform 1 0 4288 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2562
timestamp 1018054153
transform 1 0 4304 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2564
timestamp 1018054153
transform 1 0 4320 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2566
timestamp 1018054153
transform 1 0 4336 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2568
timestamp 1018054153
transform 1 0 4352 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2570
timestamp 1018054153
transform 1 0 4368 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2572
timestamp 1018054153
transform 1 0 4384 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2574
timestamp 1018054153
transform 1 0 4400 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2576
timestamp 1018054153
transform 1 0 4416 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2578
timestamp 1018054153
transform 1 0 4432 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2580
timestamp 1018054153
transform 1 0 4448 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2582
timestamp 1018054153
transform 1 0 4464 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2584
timestamp 1018054153
transform 1 0 4480 0 -1 6080
box -16 -6 32 210
use NAND2X1  NAND2X1_6
timestamp 1053022145
transform 1 0 4496 0 -1 6080
box -16 -6 64 210
use FILL  FILL_2589
timestamp 1018054153
transform 1 0 4544 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2591
timestamp 1018054153
transform 1 0 4560 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2593
timestamp 1018054153
transform 1 0 4576 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2595
timestamp 1018054153
transform 1 0 4592 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2597
timestamp 1018054153
transform 1 0 4608 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2599
timestamp 1018054153
transform 1 0 4624 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2601
timestamp 1018054153
transform 1 0 4640 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2603
timestamp 1018054153
transform 1 0 4656 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2605
timestamp 1018054153
transform 1 0 4672 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2607
timestamp 1018054153
transform 1 0 4688 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2609
timestamp 1018054153
transform 1 0 4704 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2611
timestamp 1018054153
transform 1 0 4720 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2612
timestamp 1018054153
transform 1 0 4736 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2613
timestamp 1018054153
transform 1 0 4752 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2614
timestamp 1018054153
transform 1 0 4768 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2615
timestamp 1018054153
transform 1 0 4784 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2616
timestamp 1018054153
transform 1 0 4800 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2617
timestamp 1018054153
transform 1 0 4816 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2618
timestamp 1018054153
transform 1 0 4832 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2619
timestamp 1018054153
transform 1 0 4848 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2620
timestamp 1018054153
transform 1 0 4864 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2621
timestamp 1018054153
transform 1 0 4880 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2622
timestamp 1018054153
transform 1 0 4896 0 -1 6080
box -16 -6 32 210
use NOR2X1  NOR2X1_3
timestamp 1053022145
transform 1 0 4912 0 -1 6080
box -16 -6 64 210
use FILL  FILL_2623
timestamp 1018054153
transform 1 0 4960 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2625
timestamp 1018054153
transform 1 0 4976 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2627
timestamp 1018054153
transform 1 0 4992 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2629
timestamp 1018054153
transform 1 0 5008 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2631
timestamp 1018054153
transform 1 0 5024 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2633
timestamp 1018054153
transform 1 0 5040 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2635
timestamp 1018054153
transform 1 0 5056 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2637
timestamp 1018054153
transform 1 0 5072 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2639
timestamp 1018054153
transform 1 0 5088 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2641
timestamp 1018054153
transform 1 0 5104 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2643
timestamp 1018054153
transform 1 0 5120 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2645
timestamp 1018054153
transform 1 0 5136 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2647
timestamp 1018054153
transform 1 0 5152 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2648
timestamp 1018054153
transform 1 0 5168 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2649
timestamp 1018054153
transform 1 0 5184 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2650
timestamp 1018054153
transform 1 0 5200 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2651
timestamp 1018054153
transform 1 0 5216 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2652
timestamp 1018054153
transform 1 0 5232 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2653
timestamp 1018054153
transform 1 0 5248 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2654
timestamp 1018054153
transform 1 0 5264 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2655
timestamp 1018054153
transform 1 0 5280 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2656
timestamp 1018054153
transform 1 0 5296 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2657
timestamp 1018054153
transform 1 0 5312 0 -1 6080
box -16 -6 32 210
use NOR2X1  NOR2X1_4
timestamp 1053022145
transform -1 0 5376 0 -1 6080
box -16 -6 64 210
use FILL  FILL_2658
timestamp 1018054153
transform 1 0 5376 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2659
timestamp 1018054153
transform 1 0 5392 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2661
timestamp 1018054153
transform 1 0 5408 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2663
timestamp 1018054153
transform 1 0 5424 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2665
timestamp 1018054153
transform 1 0 5440 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2667
timestamp 1018054153
transform 1 0 5456 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2669
timestamp 1018054153
transform 1 0 5472 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2671
timestamp 1018054153
transform 1 0 5488 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2673
timestamp 1018054153
transform 1 0 5504 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2675
timestamp 1018054153
transform 1 0 5520 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2677
timestamp 1018054153
transform 1 0 5536 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2679
timestamp 1018054153
transform 1 0 5552 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2681
timestamp 1018054153
transform 1 0 5568 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2683
timestamp 1018054153
transform 1 0 5584 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2685
timestamp 1018054153
transform 1 0 5600 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2693
timestamp 1018054153
transform 1 0 5616 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2694
timestamp 1018054153
transform 1 0 5632 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2695
timestamp 1018054153
transform 1 0 5648 0 -1 6080
box -16 -6 32 210
use XOR2X1  XOR2X1_1
timestamp 1053359338
transform 1 0 5664 0 -1 6080
box -16 -6 128 210
use FILL  FILL_2696
timestamp 1018054153
transform 1 0 5776 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2698
timestamp 1018054153
transform 1 0 5792 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2700
timestamp 1018054153
transform 1 0 5808 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2702
timestamp 1018054153
transform 1 0 5824 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2704
timestamp 1018054153
transform 1 0 5840 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2706
timestamp 1018054153
transform 1 0 5856 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2708
timestamp 1018054153
transform 1 0 5872 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2710
timestamp 1018054153
transform 1 0 5888 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2712
timestamp 1018054153
transform 1 0 5904 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2714
timestamp 1018054153
transform 1 0 5920 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2716
timestamp 1018054153
transform 1 0 5936 0 -1 6080
box -16 -6 32 210
use NAND3X1  NAND3X1_0
timestamp 1053022145
transform 1 0 5952 0 -1 6080
box -16 -6 80 210
use FILL  FILL_2722
timestamp 1018054153
transform 1 0 6016 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2724
timestamp 1018054153
transform 1 0 6032 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2726
timestamp 1018054153
transform 1 0 6048 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2728
timestamp 1018054153
transform 1 0 6064 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2730
timestamp 1018054153
transform 1 0 6080 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2732
timestamp 1018054153
transform 1 0 6096 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2734
timestamp 1018054153
transform 1 0 6112 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2736
timestamp 1018054153
transform 1 0 6128 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2738
timestamp 1018054153
transform 1 0 6144 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2740
timestamp 1018054153
transform 1 0 6160 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2742
timestamp 1018054153
transform 1 0 6176 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2744
timestamp 1018054153
transform 1 0 6192 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2746
timestamp 1018054153
transform 1 0 6208 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2747
timestamp 1018054153
transform 1 0 6224 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2748
timestamp 1018054153
transform 1 0 6240 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2750
timestamp 1018054153
transform 1 0 6256 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2752
timestamp 1018054153
transform 1 0 6272 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2754
timestamp 1018054153
transform 1 0 6288 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2756
timestamp 1018054153
transform 1 0 6304 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2758
timestamp 1018054153
transform 1 0 6320 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2760
timestamp 1018054153
transform 1 0 6336 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2762
timestamp 1018054153
transform 1 0 6352 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2764
timestamp 1018054153
transform 1 0 6368 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2766
timestamp 1018054153
transform 1 0 6384 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2768
timestamp 1018054153
transform 1 0 6400 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2770
timestamp 1018054153
transform 1 0 6416 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2772
timestamp 1018054153
transform 1 0 6432 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2774
timestamp 1018054153
transform 1 0 6448 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2776
timestamp 1018054153
transform 1 0 6464 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2778
timestamp 1018054153
transform 1 0 6480 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2780
timestamp 1018054153
transform 1 0 6496 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2782
timestamp 1018054153
transform 1 0 6512 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2784
timestamp 1018054153
transform 1 0 6528 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2786
timestamp 1018054153
transform 1 0 6544 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2788
timestamp 1018054153
transform 1 0 6560 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2790
timestamp 1018054153
transform 1 0 6576 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2792
timestamp 1018054153
transform 1 0 6592 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2794
timestamp 1018054153
transform 1 0 6608 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2796
timestamp 1018054153
transform 1 0 6624 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2798
timestamp 1018054153
transform 1 0 6640 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2800
timestamp 1018054153
transform 1 0 6656 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2802
timestamp 1018054153
transform 1 0 6672 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2804
timestamp 1018054153
transform 1 0 6688 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2806
timestamp 1018054153
transform 1 0 6704 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2808
timestamp 1018054153
transform 1 0 6720 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2810
timestamp 1018054153
transform 1 0 6736 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2812
timestamp 1018054153
transform 1 0 6752 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2814
timestamp 1018054153
transform 1 0 6768 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2816
timestamp 1018054153
transform 1 0 6784 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2818
timestamp 1018054153
transform 1 0 6800 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2820
timestamp 1018054153
transform 1 0 6816 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2822
timestamp 1018054153
transform 1 0 6832 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2824
timestamp 1018054153
transform 1 0 6848 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2826
timestamp 1018054153
transform 1 0 6864 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2828
timestamp 1018054153
transform 1 0 6880 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2830
timestamp 1018054153
transform 1 0 6896 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2832
timestamp 1018054153
transform 1 0 6912 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2834
timestamp 1018054153
transform 1 0 6928 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2836
timestamp 1018054153
transform 1 0 6944 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2838
timestamp 1018054153
transform 1 0 6960 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2840
timestamp 1018054153
transform 1 0 6976 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2842
timestamp 1018054153
transform 1 0 6992 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2844
timestamp 1018054153
transform 1 0 7008 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2846
timestamp 1018054153
transform 1 0 7024 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2848
timestamp 1018054153
transform 1 0 7040 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2850
timestamp 1018054153
transform 1 0 7056 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2852
timestamp 1018054153
transform 1 0 7072 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2854
timestamp 1018054153
transform 1 0 7088 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2856
timestamp 1018054153
transform 1 0 7104 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2858
timestamp 1018054153
transform 1 0 7120 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2860
timestamp 1018054153
transform 1 0 7136 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2862
timestamp 1018054153
transform 1 0 7152 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2864
timestamp 1018054153
transform 1 0 7168 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2866
timestamp 1018054153
transform 1 0 7184 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2868
timestamp 1018054153
transform 1 0 7200 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2870
timestamp 1018054153
transform 1 0 7216 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2872
timestamp 1018054153
transform 1 0 7232 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2874
timestamp 1018054153
transform 1 0 7248 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2876
timestamp 1018054153
transform 1 0 7264 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2878
timestamp 1018054153
transform 1 0 7280 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2880
timestamp 1018054153
transform 1 0 7296 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2882
timestamp 1018054153
transform 1 0 7312 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2884
timestamp 1018054153
transform 1 0 7328 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2886
timestamp 1018054153
transform 1 0 7344 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2888
timestamp 1018054153
transform 1 0 7360 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2890
timestamp 1018054153
transform 1 0 7376 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2892
timestamp 1018054153
transform 1 0 7392 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2894
timestamp 1018054153
transform 1 0 7408 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2896
timestamp 1018054153
transform 1 0 7424 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2898
timestamp 1018054153
transform 1 0 7440 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2900
timestamp 1018054153
transform 1 0 7456 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2902
timestamp 1018054153
transform 1 0 7472 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2904
timestamp 1018054153
transform 1 0 7488 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2906
timestamp 1018054153
transform 1 0 7504 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2908
timestamp 1018054153
transform 1 0 7520 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2910
timestamp 1018054153
transform 1 0 7536 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2912
timestamp 1018054153
transform 1 0 7552 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2914
timestamp 1018054153
transform 1 0 7568 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2916
timestamp 1018054153
transform 1 0 7584 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2918
timestamp 1018054153
transform 1 0 7600 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2920
timestamp 1018054153
transform 1 0 7616 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2922
timestamp 1018054153
transform 1 0 7632 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2924
timestamp 1018054153
transform 1 0 7648 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2926
timestamp 1018054153
transform 1 0 7664 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2928
timestamp 1018054153
transform 1 0 7680 0 -1 6080
box -16 -6 32 210
use FILL  FILL_2930
timestamp 1018054153
transform 1 0 7696 0 -1 6080
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_15
timestamp 1542725905
transform 1 0 7788 0 1 5880
box -48 -6 48 6
use FILL  FILL_2932
timestamp 1018054153
transform 1 0 7712 0 -1 6080
box -16 -6 32 210
use M2_M1  M2_M1_117
timestamp 1542725905
transform 1 0 3464 0 1 5750
box -4 -4 4 4
use M2_M1  M2_M1_104
timestamp 1542725905
transform 1 0 3544 0 1 5790
box -4 -4 4 4
use M2_M1  M2_M1_107
timestamp 1542725905
transform 1 0 3528 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_118
timestamp 1542725905
transform 1 0 3848 0 1 5750
box -4 -4 4 4
use M2_M1  M2_M1_105
timestamp 1542725905
transform 1 0 3912 0 1 5790
box -4 -4 4 4
use M2_M1  M2_M1_119
timestamp 1542725905
transform 1 0 4216 0 1 5750
box -4 -4 4 4
use M3_M2  M3_M2_41
timestamp 1542725905
transform 1 0 4200 0 1 5730
box -6 -6 6 6
use M2_M1  M2_M1_108
timestamp 1542725905
transform 1 0 4408 0 1 5770
box -4 -4 4 4
use M3_M2  M3_M2_37
timestamp 1542725905
transform 1 0 4440 0 1 5830
box -6 -6 6 6
use M2_M1  M2_M1_125
timestamp 1542725905
transform 1 0 4472 0 1 5730
box -4 -4 4 4
use M2_M1  M2_M1_109
timestamp 1542725905
transform 1 0 4584 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_126
timestamp 1542725905
transform 1 0 4664 0 1 5730
box -4 -4 4 4
use M2_M1  M2_M1_110
timestamp 1542725905
transform 1 0 4808 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_120
timestamp 1542725905
transform 1 0 4968 0 1 5750
box -4 -4 4 4
use M3_M2  M3_M2_39
timestamp 1542725905
transform 1 0 5112 0 1 5790
box -6 -6 6 6
use M2_M1  M2_M1_111
timestamp 1542725905
transform 1 0 5064 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_112
timestamp 1542725905
transform 1 0 5112 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_121
timestamp 1542725905
transform 1 0 5160 0 1 5750
box -4 -4 4 4
use M2_M1  M2_M1_122
timestamp 1542725905
transform 1 0 5192 0 1 5750
box -4 -4 4 4
use M3_M2  M3_M2_42
timestamp 1542725905
transform 1 0 5192 0 1 5730
box -6 -6 6 6
use M3_M2  M3_M2_40
timestamp 1542725905
transform 1 0 5224 0 1 5790
box -6 -6 6 6
use M3_M2  M3_M2_38
timestamp 1542725905
transform 1 0 5256 0 1 5830
box -6 -6 6 6
use M2_M1  M2_M1_113
timestamp 1542725905
transform 1 0 5400 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_114
timestamp 1542725905
transform 1 0 5416 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_127
timestamp 1542725905
transform 1 0 5592 0 1 5730
box -4 -4 4 4
use M2_M1  M2_M1_129
timestamp 1542725905
transform 1 0 5624 0 1 5710
box -4 -4 4 4
use M2_M1  M2_M1_130
timestamp 1542725905
transform 1 0 5720 0 1 5710
box -4 -4 4 4
use M2_M1  M2_M1_123
timestamp 1542725905
transform 1 0 5800 0 1 5750
box -4 -4 4 4
use M3_M2  M3_M2_43
timestamp 1542725905
transform 1 0 5800 0 1 5730
box -6 -6 6 6
use M2_M1  M2_M1_115
timestamp 1542725905
transform 1 0 5880 0 1 5770
box -4 -4 4 4
use M2_M1  M2_M1_106
timestamp 1542725905
transform 1 0 6024 0 1 5790
box -4 -4 4 4
use M2_M1  M2_M1_128
timestamp 1542725905
transform 1 0 6456 0 1 5730
box -4 -4 4 4
use M2_M1  M2_M1_116
timestamp 1542725905
transform 1 0 6504 0 1 5770
box -4 -4 4 4
use M3_M2  M3_M2_44
timestamp 1542725905
transform 1 0 6504 0 1 5730
box -6 -6 6 6
use M2_M1  M2_M1_124
timestamp 1542725905
transform 1 0 6568 0 1 5750
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_16
timestamp 1542725905
transform 1 0 2092 0 1 5680
box -48 -6 48 6
use FILL  FILL_2933
timestamp 1018054153
transform 1 0 2272 0 1 5680
box -16 -6 32 210
use FILL  FILL_2935
timestamp 1018054153
transform 1 0 2288 0 1 5680
box -16 -6 32 210
use FILL  FILL_2937
timestamp 1018054153
transform 1 0 2304 0 1 5680
box -16 -6 32 210
use FILL  FILL_2939
timestamp 1018054153
transform 1 0 2320 0 1 5680
box -16 -6 32 210
use FILL  FILL_2941
timestamp 1018054153
transform 1 0 2336 0 1 5680
box -16 -6 32 210
use FILL  FILL_2943
timestamp 1018054153
transform 1 0 2352 0 1 5680
box -16 -6 32 210
use FILL  FILL_2945
timestamp 1018054153
transform 1 0 2368 0 1 5680
box -16 -6 32 210
use FILL  FILL_2947
timestamp 1018054153
transform 1 0 2384 0 1 5680
box -16 -6 32 210
use FILL  FILL_2949
timestamp 1018054153
transform 1 0 2400 0 1 5680
box -16 -6 32 210
use FILL  FILL_2951
timestamp 1018054153
transform 1 0 2416 0 1 5680
box -16 -6 32 210
use FILL  FILL_2953
timestamp 1018054153
transform 1 0 2432 0 1 5680
box -16 -6 32 210
use FILL  FILL_2955
timestamp 1018054153
transform 1 0 2448 0 1 5680
box -16 -6 32 210
use FILL  FILL_2957
timestamp 1018054153
transform 1 0 2464 0 1 5680
box -16 -6 32 210
use FILL  FILL_2959
timestamp 1018054153
transform 1 0 2480 0 1 5680
box -16 -6 32 210
use FILL  FILL_2961
timestamp 1018054153
transform 1 0 2496 0 1 5680
box -16 -6 32 210
use FILL  FILL_2963
timestamp 1018054153
transform 1 0 2512 0 1 5680
box -16 -6 32 210
use FILL  FILL_2965
timestamp 1018054153
transform 1 0 2528 0 1 5680
box -16 -6 32 210
use FILL  FILL_2967
timestamp 1018054153
transform 1 0 2544 0 1 5680
box -16 -6 32 210
use FILL  FILL_2969
timestamp 1018054153
transform 1 0 2560 0 1 5680
box -16 -6 32 210
use FILL  FILL_2971
timestamp 1018054153
transform 1 0 2576 0 1 5680
box -16 -6 32 210
use FILL  FILL_2973
timestamp 1018054153
transform 1 0 2592 0 1 5680
box -16 -6 32 210
use FILL  FILL_2975
timestamp 1018054153
transform 1 0 2608 0 1 5680
box -16 -6 32 210
use FILL  FILL_2977
timestamp 1018054153
transform 1 0 2624 0 1 5680
box -16 -6 32 210
use FILL  FILL_2979
timestamp 1018054153
transform 1 0 2640 0 1 5680
box -16 -6 32 210
use FILL  FILL_2981
timestamp 1018054153
transform 1 0 2656 0 1 5680
box -16 -6 32 210
use FILL  FILL_2983
timestamp 1018054153
transform 1 0 2672 0 1 5680
box -16 -6 32 210
use FILL  FILL_2985
timestamp 1018054153
transform 1 0 2688 0 1 5680
box -16 -6 32 210
use FILL  FILL_2987
timestamp 1018054153
transform 1 0 2704 0 1 5680
box -16 -6 32 210
use FILL  FILL_2989
timestamp 1018054153
transform 1 0 2720 0 1 5680
box -16 -6 32 210
use FILL  FILL_2991
timestamp 1018054153
transform 1 0 2736 0 1 5680
box -16 -6 32 210
use FILL  FILL_2993
timestamp 1018054153
transform 1 0 2752 0 1 5680
box -16 -6 32 210
use FILL  FILL_2995
timestamp 1018054153
transform 1 0 2768 0 1 5680
box -16 -6 32 210
use FILL  FILL_2997
timestamp 1018054153
transform 1 0 2784 0 1 5680
box -16 -6 32 210
use FILL  FILL_2999
timestamp 1018054153
transform 1 0 2800 0 1 5680
box -16 -6 32 210
use FILL  FILL_3001
timestamp 1018054153
transform 1 0 2816 0 1 5680
box -16 -6 32 210
use FILL  FILL_3003
timestamp 1018054153
transform 1 0 2832 0 1 5680
box -16 -6 32 210
use FILL  FILL_3005
timestamp 1018054153
transform 1 0 2848 0 1 5680
box -16 -6 32 210
use FILL  FILL_3007
timestamp 1018054153
transform 1 0 2864 0 1 5680
box -16 -6 32 210
use FILL  FILL_3009
timestamp 1018054153
transform 1 0 2880 0 1 5680
box -16 -6 32 210
use FILL  FILL_3011
timestamp 1018054153
transform 1 0 2896 0 1 5680
box -16 -6 32 210
use FILL  FILL_3013
timestamp 1018054153
transform 1 0 2912 0 1 5680
box -16 -6 32 210
use FILL  FILL_3015
timestamp 1018054153
transform 1 0 2928 0 1 5680
box -16 -6 32 210
use FILL  FILL_3017
timestamp 1018054153
transform 1 0 2944 0 1 5680
box -16 -6 32 210
use FILL  FILL_3019
timestamp 1018054153
transform 1 0 2960 0 1 5680
box -16 -6 32 210
use FILL  FILL_3021
timestamp 1018054153
transform 1 0 2976 0 1 5680
box -16 -6 32 210
use FILL  FILL_3023
timestamp 1018054153
transform 1 0 2992 0 1 5680
box -16 -6 32 210
use FILL  FILL_3025
timestamp 1018054153
transform 1 0 3008 0 1 5680
box -16 -6 32 210
use FILL  FILL_3027
timestamp 1018054153
transform 1 0 3024 0 1 5680
box -16 -6 32 210
use FILL  FILL_3029
timestamp 1018054153
transform 1 0 3040 0 1 5680
box -16 -6 32 210
use FILL  FILL_3031
timestamp 1018054153
transform 1 0 3056 0 1 5680
box -16 -6 32 210
use FILL  FILL_3033
timestamp 1018054153
transform 1 0 3072 0 1 5680
box -16 -6 32 210
use FILL  FILL_3035
timestamp 1018054153
transform 1 0 3088 0 1 5680
box -16 -6 32 210
use FILL  FILL_3037
timestamp 1018054153
transform 1 0 3104 0 1 5680
box -16 -6 32 210
use FILL  FILL_3039
timestamp 1018054153
transform 1 0 3120 0 1 5680
box -16 -6 32 210
use FILL  FILL_3041
timestamp 1018054153
transform 1 0 3136 0 1 5680
box -16 -6 32 210
use FILL  FILL_3043
timestamp 1018054153
transform 1 0 3152 0 1 5680
box -16 -6 32 210
use FILL  FILL_3045
timestamp 1018054153
transform 1 0 3168 0 1 5680
box -16 -6 32 210
use FILL  FILL_3047
timestamp 1018054153
transform 1 0 3184 0 1 5680
box -16 -6 32 210
use FILL  FILL_3049
timestamp 1018054153
transform 1 0 3200 0 1 5680
box -16 -6 32 210
use FILL  FILL_3051
timestamp 1018054153
transform 1 0 3216 0 1 5680
box -16 -6 32 210
use FILL  FILL_3053
timestamp 1018054153
transform 1 0 3232 0 1 5680
box -16 -6 32 210
use FILL  FILL_3055
timestamp 1018054153
transform 1 0 3248 0 1 5680
box -16 -6 32 210
use FILL  FILL_3057
timestamp 1018054153
transform 1 0 3264 0 1 5680
box -16 -6 32 210
use FILL  FILL_3059
timestamp 1018054153
transform 1 0 3280 0 1 5680
box -16 -6 32 210
use FILL  FILL_3061
timestamp 1018054153
transform 1 0 3296 0 1 5680
box -16 -6 32 210
use FILL  FILL_3063
timestamp 1018054153
transform 1 0 3312 0 1 5680
box -16 -6 32 210
use FILL  FILL_3065
timestamp 1018054153
transform 1 0 3328 0 1 5680
box -16 -6 32 210
use FILL  FILL_3067
timestamp 1018054153
transform 1 0 3344 0 1 5680
box -16 -6 32 210
use FILL  FILL_3069
timestamp 1018054153
transform 1 0 3360 0 1 5680
box -16 -6 32 210
use FILL  FILL_3071
timestamp 1018054153
transform 1 0 3376 0 1 5680
box -16 -6 32 210
use FILL  FILL_3073
timestamp 1018054153
transform 1 0 3392 0 1 5680
box -16 -6 32 210
use FILL  FILL_3075
timestamp 1018054153
transform 1 0 3408 0 1 5680
box -16 -6 32 210
use FILL  FILL_3077
timestamp 1018054153
transform 1 0 3424 0 1 5680
box -16 -6 32 210
use FILL  FILL_3079
timestamp 1018054153
transform 1 0 3440 0 1 5680
box -16 -6 32 210
use FILL  FILL_3081
timestamp 1018054153
transform 1 0 3456 0 1 5680
box -16 -6 32 210
use FILL  FILL_3083
timestamp 1018054153
transform 1 0 3472 0 1 5680
box -16 -6 32 210
use FILL  FILL_3085
timestamp 1018054153
transform 1 0 3488 0 1 5680
box -16 -6 32 210
use NAND2X1  NAND2X1_7
timestamp 1053022145
transform 1 0 3504 0 1 5680
box -16 -6 64 210
use FILL  FILL_3087
timestamp 1018054153
transform 1 0 3552 0 1 5680
box -16 -6 32 210
use FILL  FILL_3092
timestamp 1018054153
transform 1 0 3568 0 1 5680
box -16 -6 32 210
use FILL  FILL_3094
timestamp 1018054153
transform 1 0 3584 0 1 5680
box -16 -6 32 210
use FILL  FILL_3096
timestamp 1018054153
transform 1 0 3600 0 1 5680
box -16 -6 32 210
use FILL  FILL_3098
timestamp 1018054153
transform 1 0 3616 0 1 5680
box -16 -6 32 210
use FILL  FILL_3100
timestamp 1018054153
transform 1 0 3632 0 1 5680
box -16 -6 32 210
use FILL  FILL_3102
timestamp 1018054153
transform 1 0 3648 0 1 5680
box -16 -6 32 210
use FILL  FILL_3104
timestamp 1018054153
transform 1 0 3664 0 1 5680
box -16 -6 32 210
use FILL  FILL_3106
timestamp 1018054153
transform 1 0 3680 0 1 5680
box -16 -6 32 210
use FILL  FILL_3108
timestamp 1018054153
transform 1 0 3696 0 1 5680
box -16 -6 32 210
use FILL  FILL_3110
timestamp 1018054153
transform 1 0 3712 0 1 5680
box -16 -6 32 210
use FILL  FILL_3112
timestamp 1018054153
transform 1 0 3728 0 1 5680
box -16 -6 32 210
use FILL  FILL_3114
timestamp 1018054153
transform 1 0 3744 0 1 5680
box -16 -6 32 210
use FILL  FILL_3116
timestamp 1018054153
transform 1 0 3760 0 1 5680
box -16 -6 32 210
use FILL  FILL_3118
timestamp 1018054153
transform 1 0 3776 0 1 5680
box -16 -6 32 210
use FILL  FILL_3120
timestamp 1018054153
transform 1 0 3792 0 1 5680
box -16 -6 32 210
use FILL  FILL_3122
timestamp 1018054153
transform 1 0 3808 0 1 5680
box -16 -6 32 210
use FILL  FILL_3124
timestamp 1018054153
transform 1 0 3824 0 1 5680
box -16 -6 32 210
use FILL  FILL_3126
timestamp 1018054153
transform 1 0 3840 0 1 5680
box -16 -6 32 210
use FILL  FILL_3127
timestamp 1018054153
transform 1 0 3856 0 1 5680
box -16 -6 32 210
use FILL  FILL_3128
timestamp 1018054153
transform 1 0 3872 0 1 5680
box -16 -6 32 210
use FILL  FILL_3129
timestamp 1018054153
transform 1 0 3888 0 1 5680
box -16 -6 32 210
use FILL  FILL_3130
timestamp 1018054153
transform 1 0 3904 0 1 5680
box -16 -6 32 210
use FILL  FILL_3132
timestamp 1018054153
transform 1 0 3920 0 1 5680
box -16 -6 32 210
use FILL  FILL_3134
timestamp 1018054153
transform 1 0 3936 0 1 5680
box -16 -6 32 210
use FILL  FILL_3136
timestamp 1018054153
transform 1 0 3952 0 1 5680
box -16 -6 32 210
use FILL  FILL_3138
timestamp 1018054153
transform 1 0 3968 0 1 5680
box -16 -6 32 210
use FILL  FILL_3140
timestamp 1018054153
transform 1 0 3984 0 1 5680
box -16 -6 32 210
use FILL  FILL_3142
timestamp 1018054153
transform 1 0 4000 0 1 5680
box -16 -6 32 210
use FILL  FILL_3144
timestamp 1018054153
transform 1 0 4016 0 1 5680
box -16 -6 32 210
use M3_M2  M3_M2_45
timestamp 1542725905
transform 1 0 4056 0 1 5690
box -6 -6 6 6
use FILL  FILL_3146
timestamp 1018054153
transform 1 0 4032 0 1 5680
box -16 -6 32 210
use FILL  FILL_3148
timestamp 1018054153
transform 1 0 4048 0 1 5680
box -16 -6 32 210
use FILL  FILL_3150
timestamp 1018054153
transform 1 0 4064 0 1 5680
box -16 -6 32 210
use FILL  FILL_3152
timestamp 1018054153
transform 1 0 4080 0 1 5680
box -16 -6 32 210
use FILL  FILL_3154
timestamp 1018054153
transform 1 0 4096 0 1 5680
box -16 -6 32 210
use FILL  FILL_3156
timestamp 1018054153
transform 1 0 4112 0 1 5680
box -16 -6 32 210
use FILL  FILL_3158
timestamp 1018054153
transform 1 0 4128 0 1 5680
box -16 -6 32 210
use FILL  FILL_3160
timestamp 1018054153
transform 1 0 4144 0 1 5680
box -16 -6 32 210
use FILL  FILL_3162
timestamp 1018054153
transform 1 0 4160 0 1 5680
box -16 -6 32 210
use FILL  FILL_3164
timestamp 1018054153
transform 1 0 4176 0 1 5680
box -16 -6 32 210
use FILL  FILL_3166
timestamp 1018054153
transform 1 0 4192 0 1 5680
box -16 -6 32 210
use FILL  FILL_3168
timestamp 1018054153
transform 1 0 4208 0 1 5680
box -16 -6 32 210
use FILL  FILL_3170
timestamp 1018054153
transform 1 0 4224 0 1 5680
box -16 -6 32 210
use FILL  FILL_3172
timestamp 1018054153
transform 1 0 4240 0 1 5680
box -16 -6 32 210
use FILL  FILL_3174
timestamp 1018054153
transform 1 0 4256 0 1 5680
box -16 -6 32 210
use FILL  FILL_3176
timestamp 1018054153
transform 1 0 4272 0 1 5680
box -16 -6 32 210
use FILL  FILL_3178
timestamp 1018054153
transform 1 0 4288 0 1 5680
box -16 -6 32 210
use FILL  FILL_3180
timestamp 1018054153
transform 1 0 4304 0 1 5680
box -16 -6 32 210
use FILL  FILL_3182
timestamp 1018054153
transform 1 0 4320 0 1 5680
box -16 -6 32 210
use FILL  FILL_3184
timestamp 1018054153
transform 1 0 4336 0 1 5680
box -16 -6 32 210
use FILL  FILL_3186
timestamp 1018054153
transform 1 0 4352 0 1 5680
box -16 -6 32 210
use FILL  FILL_3188
timestamp 1018054153
transform 1 0 4368 0 1 5680
box -16 -6 32 210
use FILL  FILL_3190
timestamp 1018054153
transform 1 0 4384 0 1 5680
box -16 -6 32 210
use FILL  FILL_3192
timestamp 1018054153
transform 1 0 4400 0 1 5680
box -16 -6 32 210
use AOI21X1  AOI21X1_1
timestamp 1090541997
transform 1 0 4416 0 1 5680
box -14 -6 78 210
use FILL  FILL_3194
timestamp 1018054153
transform 1 0 4480 0 1 5680
box -16 -6 32 210
use FILL  FILL_3195
timestamp 1018054153
transform 1 0 4496 0 1 5680
box -16 -6 32 210
use FILL  FILL_3197
timestamp 1018054153
transform 1 0 4512 0 1 5680
box -16 -6 32 210
use FILL  FILL_3199
timestamp 1018054153
transform 1 0 4528 0 1 5680
box -16 -6 32 210
use FILL  FILL_3201
timestamp 1018054153
transform 1 0 4544 0 1 5680
box -16 -6 32 210
use FILL  FILL_3203
timestamp 1018054153
transform 1 0 4560 0 1 5680
box -16 -6 32 210
use FILL  FILL_3205
timestamp 1018054153
transform 1 0 4576 0 1 5680
box -16 -6 32 210
use FILL  FILL_3207
timestamp 1018054153
transform 1 0 4592 0 1 5680
box -16 -6 32 210
use FILL  FILL_3209
timestamp 1018054153
transform 1 0 4608 0 1 5680
box -16 -6 32 210
use FILL  FILL_3211
timestamp 1018054153
transform 1 0 4624 0 1 5680
box -16 -6 32 210
use M3_M2  M3_M2_46
timestamp 1542725905
transform 1 0 4664 0 1 5690
box -6 -6 6 6
use FILL  FILL_3213
timestamp 1018054153
transform 1 0 4640 0 1 5680
box -16 -6 32 210
use FILL  FILL_3215
timestamp 1018054153
transform 1 0 4656 0 1 5680
box -16 -6 32 210
use FILL  FILL_3217
timestamp 1018054153
transform 1 0 4672 0 1 5680
box -16 -6 32 210
use FILL  FILL_3219
timestamp 1018054153
transform 1 0 4688 0 1 5680
box -16 -6 32 210
use FILL  FILL_3221
timestamp 1018054153
transform 1 0 4704 0 1 5680
box -16 -6 32 210
use FILL  FILL_3223
timestamp 1018054153
transform 1 0 4720 0 1 5680
box -16 -6 32 210
use FILL  FILL_3225
timestamp 1018054153
transform 1 0 4736 0 1 5680
box -16 -6 32 210
use FILL  FILL_3227
timestamp 1018054153
transform 1 0 4752 0 1 5680
box -16 -6 32 210
use NOR2X1  NOR2X1_5
timestamp 1053022145
transform 1 0 4768 0 1 5680
box -16 -6 64 210
use FILL  FILL_3229
timestamp 1018054153
transform 1 0 4816 0 1 5680
box -16 -6 32 210
use FILL  FILL_3234
timestamp 1018054153
transform 1 0 4832 0 1 5680
box -16 -6 32 210
use FILL  FILL_3236
timestamp 1018054153
transform 1 0 4848 0 1 5680
box -16 -6 32 210
use FILL  FILL_3238
timestamp 1018054153
transform 1 0 4864 0 1 5680
box -16 -6 32 210
use FILL  FILL_3240
timestamp 1018054153
transform 1 0 4880 0 1 5680
box -16 -6 32 210
use FILL  FILL_3242
timestamp 1018054153
transform 1 0 4896 0 1 5680
box -16 -6 32 210
use FILL  FILL_3243
timestamp 1018054153
transform 1 0 4912 0 1 5680
box -16 -6 32 210
use FILL  FILL_3244
timestamp 1018054153
transform 1 0 4928 0 1 5680
box -16 -6 32 210
use FILL  FILL_3245
timestamp 1018054153
transform 1 0 4944 0 1 5680
box -16 -6 32 210
use FILL  FILL_3248
timestamp 1018054153
transform 1 0 4960 0 1 5680
box -16 -6 32 210
use FILL  FILL_3250
timestamp 1018054153
transform 1 0 4976 0 1 5680
box -16 -6 32 210
use FILL  FILL_3252
timestamp 1018054153
transform 1 0 4992 0 1 5680
box -16 -6 32 210
use FILL  FILL_3254
timestamp 1018054153
transform 1 0 5008 0 1 5680
box -16 -6 32 210
use FILL  FILL_3256
timestamp 1018054153
transform 1 0 5024 0 1 5680
box -16 -6 32 210
use FILL  FILL_3258
timestamp 1018054153
transform 1 0 5040 0 1 5680
box -16 -6 32 210
use XOR2X1  XOR2X1_2
timestamp 1053359338
transform -1 0 5168 0 1 5680
box -16 -6 128 210
use FILL  FILL_3259
timestamp 1018054153
transform 1 0 5168 0 1 5680
box -16 -6 32 210
use FILL  FILL_3269
timestamp 1018054153
transform 1 0 5184 0 1 5680
box -16 -6 32 210
use FILL  FILL_3270
timestamp 1018054153
transform 1 0 5200 0 1 5680
box -16 -6 32 210
use FILL  FILL_3271
timestamp 1018054153
transform 1 0 5216 0 1 5680
box -16 -6 32 210
use FILL  FILL_3272
timestamp 1018054153
transform 1 0 5232 0 1 5680
box -16 -6 32 210
use FILL  FILL_3274
timestamp 1018054153
transform 1 0 5248 0 1 5680
box -16 -6 32 210
use FILL  FILL_3276
timestamp 1018054153
transform 1 0 5264 0 1 5680
box -16 -6 32 210
use FILL  FILL_3278
timestamp 1018054153
transform 1 0 5280 0 1 5680
box -16 -6 32 210
use FILL  FILL_3280
timestamp 1018054153
transform 1 0 5296 0 1 5680
box -16 -6 32 210
use FILL  FILL_3282
timestamp 1018054153
transform 1 0 5312 0 1 5680
box -16 -6 32 210
use FILL  FILL_3284
timestamp 1018054153
transform 1 0 5328 0 1 5680
box -16 -6 32 210
use FILL  FILL_3286
timestamp 1018054153
transform 1 0 5344 0 1 5680
box -16 -6 32 210
use FILL  FILL_3288
timestamp 1018054153
transform 1 0 5360 0 1 5680
box -16 -6 32 210
use FAX1  FAX1_2
timestamp 1053025068
transform 1 0 5376 0 1 5680
box -10 -6 252 210
use FILL  FILL_3290
timestamp 1018054153
transform 1 0 5616 0 1 5680
box -16 -6 32 210
use FILL  FILL_3304
timestamp 1018054153
transform 1 0 5632 0 1 5680
box -16 -6 32 210
use FILL  FILL_3306
timestamp 1018054153
transform 1 0 5648 0 1 5680
box -16 -6 32 210
use FILL  FILL_3308
timestamp 1018054153
transform 1 0 5664 0 1 5680
box -16 -6 32 210
use FILL  FILL_3310
timestamp 1018054153
transform 1 0 5680 0 1 5680
box -16 -6 32 210
use FILL  FILL_3312
timestamp 1018054153
transform 1 0 5696 0 1 5680
box -16 -6 32 210
use FILL  FILL_3314
timestamp 1018054153
transform 1 0 5712 0 1 5680
box -16 -6 32 210
use FILL  FILL_3316
timestamp 1018054153
transform 1 0 5728 0 1 5680
box -16 -6 32 210
use FILL  FILL_3318
timestamp 1018054153
transform 1 0 5744 0 1 5680
box -16 -6 32 210
use FILL  FILL_3320
timestamp 1018054153
transform 1 0 5760 0 1 5680
box -16 -6 32 210
use FILL  FILL_3322
timestamp 1018054153
transform 1 0 5776 0 1 5680
box -16 -6 32 210
use FILL  FILL_3324
timestamp 1018054153
transform 1 0 5792 0 1 5680
box -16 -6 32 210
use FILL  FILL_3326
timestamp 1018054153
transform 1 0 5808 0 1 5680
box -16 -6 32 210
use FILL  FILL_3328
timestamp 1018054153
transform 1 0 5824 0 1 5680
box -16 -6 32 210
use FILL  FILL_3330
timestamp 1018054153
transform 1 0 5840 0 1 5680
box -16 -6 32 210
use OAI21X1  OAI21X1_10
timestamp 1053722159
transform 1 0 5856 0 1 5680
box -16 -6 68 210
use FILL  FILL_3332
timestamp 1018054153
transform 1 0 5920 0 1 5680
box -16 -6 32 210
use FILL  FILL_3333
timestamp 1018054153
transform 1 0 5936 0 1 5680
box -16 -6 32 210
use FILL  FILL_3334
timestamp 1018054153
transform 1 0 5952 0 1 5680
box -16 -6 32 210
use FILL  FILL_3335
timestamp 1018054153
transform 1 0 5968 0 1 5680
box -16 -6 32 210
use FILL  FILL_3336
timestamp 1018054153
transform 1 0 5984 0 1 5680
box -16 -6 32 210
use FILL  FILL_3343
timestamp 1018054153
transform 1 0 6000 0 1 5680
box -16 -6 32 210
use FILL  FILL_3345
timestamp 1018054153
transform 1 0 6016 0 1 5680
box -16 -6 32 210
use FILL  FILL_3347
timestamp 1018054153
transform 1 0 6032 0 1 5680
box -16 -6 32 210
use FILL  FILL_3349
timestamp 1018054153
transform 1 0 6048 0 1 5680
box -16 -6 32 210
use FILL  FILL_3351
timestamp 1018054153
transform 1 0 6064 0 1 5680
box -16 -6 32 210
use FILL  FILL_3353
timestamp 1018054153
transform 1 0 6080 0 1 5680
box -16 -6 32 210
use FILL  FILL_3355
timestamp 1018054153
transform 1 0 6096 0 1 5680
box -16 -6 32 210
use FILL  FILL_3357
timestamp 1018054153
transform 1 0 6112 0 1 5680
box -16 -6 32 210
use FILL  FILL_3359
timestamp 1018054153
transform 1 0 6128 0 1 5680
box -16 -6 32 210
use FILL  FILL_3361
timestamp 1018054153
transform 1 0 6144 0 1 5680
box -16 -6 32 210
use FILL  FILL_3363
timestamp 1018054153
transform 1 0 6160 0 1 5680
box -16 -6 32 210
use FILL  FILL_3365
timestamp 1018054153
transform 1 0 6176 0 1 5680
box -16 -6 32 210
use INVX1  INVX1_7
timestamp 1053022145
transform 1 0 6192 0 1 5680
box -18 -6 52 210
use FILL  FILL_3366
timestamp 1018054153
transform 1 0 6224 0 1 5680
box -16 -6 32 210
use FILL  FILL_3369
timestamp 1018054153
transform 1 0 6240 0 1 5680
box -16 -6 32 210
use FILL  FILL_3371
timestamp 1018054153
transform 1 0 6256 0 1 5680
box -16 -6 32 210
use FILL  FILL_3373
timestamp 1018054153
transform 1 0 6272 0 1 5680
box -16 -6 32 210
use FILL  FILL_3375
timestamp 1018054153
transform 1 0 6288 0 1 5680
box -16 -6 32 210
use FILL  FILL_3377
timestamp 1018054153
transform 1 0 6304 0 1 5680
box -16 -6 32 210
use FILL  FILL_3379
timestamp 1018054153
transform 1 0 6320 0 1 5680
box -16 -6 32 210
use FILL  FILL_3381
timestamp 1018054153
transform 1 0 6336 0 1 5680
box -16 -6 32 210
use FILL  FILL_3383
timestamp 1018054153
transform 1 0 6352 0 1 5680
box -16 -6 32 210
use FILL  FILL_3385
timestamp 1018054153
transform 1 0 6368 0 1 5680
box -16 -6 32 210
use FILL  FILL_3387
timestamp 1018054153
transform 1 0 6384 0 1 5680
box -16 -6 32 210
use FILL  FILL_3389
timestamp 1018054153
transform 1 0 6400 0 1 5680
box -16 -6 32 210
use FILL  FILL_3391
timestamp 1018054153
transform 1 0 6416 0 1 5680
box -16 -6 32 210
use FILL  FILL_3393
timestamp 1018054153
transform 1 0 6432 0 1 5680
box -16 -6 32 210
use FILL  FILL_3395
timestamp 1018054153
transform 1 0 6448 0 1 5680
box -16 -6 32 210
use NOR2X1  NOR2X1_7
timestamp 1053022145
transform 1 0 6464 0 1 5680
box -16 -6 64 210
use FILL  FILL_3397
timestamp 1018054153
transform 1 0 6512 0 1 5680
box -16 -6 32 210
use FILL  FILL_3398
timestamp 1018054153
transform 1 0 6528 0 1 5680
box -16 -6 32 210
use FILL  FILL_3399
timestamp 1018054153
transform 1 0 6544 0 1 5680
box -16 -6 32 210
use FILL  FILL_3400
timestamp 1018054153
transform 1 0 6560 0 1 5680
box -16 -6 32 210
use FILL  FILL_3404
timestamp 1018054153
transform 1 0 6576 0 1 5680
box -16 -6 32 210
use FILL  FILL_3406
timestamp 1018054153
transform 1 0 6592 0 1 5680
box -16 -6 32 210
use FILL  FILL_3408
timestamp 1018054153
transform 1 0 6608 0 1 5680
box -16 -6 32 210
use FILL  FILL_3410
timestamp 1018054153
transform 1 0 6624 0 1 5680
box -16 -6 32 210
use FILL  FILL_3412
timestamp 1018054153
transform 1 0 6640 0 1 5680
box -16 -6 32 210
use FILL  FILL_3414
timestamp 1018054153
transform 1 0 6656 0 1 5680
box -16 -6 32 210
use FILL  FILL_3416
timestamp 1018054153
transform 1 0 6672 0 1 5680
box -16 -6 32 210
use FILL  FILL_3418
timestamp 1018054153
transform 1 0 6688 0 1 5680
box -16 -6 32 210
use FILL  FILL_3420
timestamp 1018054153
transform 1 0 6704 0 1 5680
box -16 -6 32 210
use FILL  FILL_3422
timestamp 1018054153
transform 1 0 6720 0 1 5680
box -16 -6 32 210
use FILL  FILL_3424
timestamp 1018054153
transform 1 0 6736 0 1 5680
box -16 -6 32 210
use FILL  FILL_3426
timestamp 1018054153
transform 1 0 6752 0 1 5680
box -16 -6 32 210
use FILL  FILL_3428
timestamp 1018054153
transform 1 0 6768 0 1 5680
box -16 -6 32 210
use FILL  FILL_3430
timestamp 1018054153
transform 1 0 6784 0 1 5680
box -16 -6 32 210
use FILL  FILL_3432
timestamp 1018054153
transform 1 0 6800 0 1 5680
box -16 -6 32 210
use FILL  FILL_3434
timestamp 1018054153
transform 1 0 6816 0 1 5680
box -16 -6 32 210
use FILL  FILL_3436
timestamp 1018054153
transform 1 0 6832 0 1 5680
box -16 -6 32 210
use FILL  FILL_3438
timestamp 1018054153
transform 1 0 6848 0 1 5680
box -16 -6 32 210
use FILL  FILL_3440
timestamp 1018054153
transform 1 0 6864 0 1 5680
box -16 -6 32 210
use FILL  FILL_3442
timestamp 1018054153
transform 1 0 6880 0 1 5680
box -16 -6 32 210
use FILL  FILL_3444
timestamp 1018054153
transform 1 0 6896 0 1 5680
box -16 -6 32 210
use FILL  FILL_3446
timestamp 1018054153
transform 1 0 6912 0 1 5680
box -16 -6 32 210
use FILL  FILL_3448
timestamp 1018054153
transform 1 0 6928 0 1 5680
box -16 -6 32 210
use FILL  FILL_3450
timestamp 1018054153
transform 1 0 6944 0 1 5680
box -16 -6 32 210
use FILL  FILL_3452
timestamp 1018054153
transform 1 0 6960 0 1 5680
box -16 -6 32 210
use FILL  FILL_3454
timestamp 1018054153
transform 1 0 6976 0 1 5680
box -16 -6 32 210
use FILL  FILL_3456
timestamp 1018054153
transform 1 0 6992 0 1 5680
box -16 -6 32 210
use FILL  FILL_3458
timestamp 1018054153
transform 1 0 7008 0 1 5680
box -16 -6 32 210
use FILL  FILL_3460
timestamp 1018054153
transform 1 0 7024 0 1 5680
box -16 -6 32 210
use FILL  FILL_3462
timestamp 1018054153
transform 1 0 7040 0 1 5680
box -16 -6 32 210
use FILL  FILL_3464
timestamp 1018054153
transform 1 0 7056 0 1 5680
box -16 -6 32 210
use FILL  FILL_3466
timestamp 1018054153
transform 1 0 7072 0 1 5680
box -16 -6 32 210
use FILL  FILL_3468
timestamp 1018054153
transform 1 0 7088 0 1 5680
box -16 -6 32 210
use FILL  FILL_3470
timestamp 1018054153
transform 1 0 7104 0 1 5680
box -16 -6 32 210
use FILL  FILL_3472
timestamp 1018054153
transform 1 0 7120 0 1 5680
box -16 -6 32 210
use FILL  FILL_3474
timestamp 1018054153
transform 1 0 7136 0 1 5680
box -16 -6 32 210
use FILL  FILL_3476
timestamp 1018054153
transform 1 0 7152 0 1 5680
box -16 -6 32 210
use FILL  FILL_3478
timestamp 1018054153
transform 1 0 7168 0 1 5680
box -16 -6 32 210
use FILL  FILL_3480
timestamp 1018054153
transform 1 0 7184 0 1 5680
box -16 -6 32 210
use FILL  FILL_3482
timestamp 1018054153
transform 1 0 7200 0 1 5680
box -16 -6 32 210
use FILL  FILL_3484
timestamp 1018054153
transform 1 0 7216 0 1 5680
box -16 -6 32 210
use FILL  FILL_3486
timestamp 1018054153
transform 1 0 7232 0 1 5680
box -16 -6 32 210
use FILL  FILL_3488
timestamp 1018054153
transform 1 0 7248 0 1 5680
box -16 -6 32 210
use FILL  FILL_3490
timestamp 1018054153
transform 1 0 7264 0 1 5680
box -16 -6 32 210
use FILL  FILL_3492
timestamp 1018054153
transform 1 0 7280 0 1 5680
box -16 -6 32 210
use FILL  FILL_3494
timestamp 1018054153
transform 1 0 7296 0 1 5680
box -16 -6 32 210
use FILL  FILL_3496
timestamp 1018054153
transform 1 0 7312 0 1 5680
box -16 -6 32 210
use FILL  FILL_3498
timestamp 1018054153
transform 1 0 7328 0 1 5680
box -16 -6 32 210
use FILL  FILL_3500
timestamp 1018054153
transform 1 0 7344 0 1 5680
box -16 -6 32 210
use FILL  FILL_3502
timestamp 1018054153
transform 1 0 7360 0 1 5680
box -16 -6 32 210
use FILL  FILL_3504
timestamp 1018054153
transform 1 0 7376 0 1 5680
box -16 -6 32 210
use FILL  FILL_3506
timestamp 1018054153
transform 1 0 7392 0 1 5680
box -16 -6 32 210
use FILL  FILL_3508
timestamp 1018054153
transform 1 0 7408 0 1 5680
box -16 -6 32 210
use FILL  FILL_3510
timestamp 1018054153
transform 1 0 7424 0 1 5680
box -16 -6 32 210
use FILL  FILL_3512
timestamp 1018054153
transform 1 0 7440 0 1 5680
box -16 -6 32 210
use FILL  FILL_3514
timestamp 1018054153
transform 1 0 7456 0 1 5680
box -16 -6 32 210
use FILL  FILL_3516
timestamp 1018054153
transform 1 0 7472 0 1 5680
box -16 -6 32 210
use FILL  FILL_3518
timestamp 1018054153
transform 1 0 7488 0 1 5680
box -16 -6 32 210
use FILL  FILL_3520
timestamp 1018054153
transform 1 0 7504 0 1 5680
box -16 -6 32 210
use FILL  FILL_3522
timestamp 1018054153
transform 1 0 7520 0 1 5680
box -16 -6 32 210
use FILL  FILL_3524
timestamp 1018054153
transform 1 0 7536 0 1 5680
box -16 -6 32 210
use FILL  FILL_3526
timestamp 1018054153
transform 1 0 7552 0 1 5680
box -16 -6 32 210
use FILL  FILL_3528
timestamp 1018054153
transform 1 0 7568 0 1 5680
box -16 -6 32 210
use FILL  FILL_3530
timestamp 1018054153
transform 1 0 7584 0 1 5680
box -16 -6 32 210
use FILL  FILL_3532
timestamp 1018054153
transform 1 0 7600 0 1 5680
box -16 -6 32 210
use FILL  FILL_3534
timestamp 1018054153
transform 1 0 7616 0 1 5680
box -16 -6 32 210
use FILL  FILL_3536
timestamp 1018054153
transform 1 0 7632 0 1 5680
box -16 -6 32 210
use FILL  FILL_3538
timestamp 1018054153
transform 1 0 7648 0 1 5680
box -16 -6 32 210
use FILL  FILL_3540
timestamp 1018054153
transform 1 0 7664 0 1 5680
box -16 -6 32 210
use FILL  FILL_3542
timestamp 1018054153
transform 1 0 7680 0 1 5680
box -16 -6 32 210
use FILL  FILL_3544
timestamp 1018054153
transform 1 0 7696 0 1 5680
box -16 -6 32 210
use FILL  FILL_3546
timestamp 1018054153
transform 1 0 7712 0 1 5680
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_17
timestamp 1542725905
transform 1 0 7908 0 1 5680
box -48 -6 48 6
use PADINC  PADINC_5
timestamp 1084294328
transform 0 -1 2000 1 0 5600
box -12 -6 606 2000
use M3_M2  M3_M2_50
timestamp 1542725905
transform 1 0 1998 0 1 5530
box -6 -6 6 6
use M3_M2  M3_M2_47
timestamp 1542725905
transform 1 0 3048 0 1 5570
box -6 -6 6 6
use M2_M1  M2_M1_148
timestamp 1542725905
transform 1 0 3464 0 1 5590
box -4 -4 4 4
use M2_M1  M2_M1_136
timestamp 1542725905
transform 1 0 3848 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_154
timestamp 1542725905
transform 1 0 3912 0 1 5570
box -4 -4 4 4
use M3_M2  M3_M2_48
timestamp 1542725905
transform 1 0 4104 0 1 5570
box -6 -6 6 6
use M2_M1  M2_M1_137
timestamp 1542725905
transform 1 0 4200 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_149
timestamp 1542725905
transform 1 0 4216 0 1 5590
box -4 -4 4 4
use M2_M1  M2_M1_138
timestamp 1542725905
transform 1 0 4440 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_139
timestamp 1542725905
transform 1 0 4472 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_150
timestamp 1542725905
transform 1 0 4456 0 1 5590
box -4 -4 4 4
use M2_M1  M2_M1_151
timestamp 1542725905
transform 1 0 4520 0 1 5590
box -4 -4 4 4
use M3_M2  M3_M2_51
timestamp 1542725905
transform 1 0 4520 0 1 5530
box -6 -6 6 6
use M2_M1  M2_M1_140
timestamp 1542725905
transform 1 0 4552 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_141
timestamp 1542725905
transform 1 0 4920 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_132
timestamp 1542725905
transform 1 0 4968 0 1 5630
box -4 -4 4 4
use M2_M1  M2_M1_133
timestamp 1542725905
transform 1 0 5048 0 1 5630
box -4 -4 4 4
use M2_M1  M2_M1_142
timestamp 1542725905
transform 1 0 5080 0 1 5610
box -4 -4 4 4
use M3_M2  M3_M2_49
timestamp 1542725905
transform 1 0 5080 0 1 5570
box -6 -6 6 6
use M2_M1  M2_M1_155
timestamp 1542725905
transform 1 0 5256 0 1 5570
box -4 -4 4 4
use M2_M1  M2_M1_134
timestamp 1542725905
transform 1 0 5416 0 1 5630
box -4 -4 4 4
use M2_M1  M2_M1_143
timestamp 1542725905
transform 1 0 5400 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_156
timestamp 1542725905
transform 1 0 5512 0 1 5570
box -4 -4 4 4
use M3_M2  M3_M2_52
timestamp 1542725905
transform 1 0 5512 0 1 5530
box -6 -6 6 6
use M2_M1  M2_M1_144
timestamp 1542725905
transform 1 0 5560 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_145
timestamp 1542725905
transform 1 0 5880 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_146
timestamp 1542725905
transform 1 0 5992 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_131
timestamp 1542725905
transform 1 0 6024 0 1 5650
box -4 -4 4 4
use M2_M1  M2_M1_147
timestamp 1542725905
transform 1 0 6472 0 1 5610
box -4 -4 4 4
use M2_M1  M2_M1_152
timestamp 1542725905
transform 1 0 6504 0 1 5590
box -4 -4 4 4
use M2_M1  M2_M1_135
timestamp 1542725905
transform 1 0 6568 0 1 5630
box -4 -4 4 4
use M2_M1  M2_M1_153
timestamp 1542725905
transform 1 0 6600 0 1 5590
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_18
timestamp 1542725905
transform 1 0 2212 0 1 5480
box -48 -6 48 6
use FILL  FILL_2934
timestamp 1018054153
transform 1 0 2272 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2936
timestamp 1018054153
transform 1 0 2288 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2938
timestamp 1018054153
transform 1 0 2304 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2940
timestamp 1018054153
transform 1 0 2320 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2942
timestamp 1018054153
transform 1 0 2336 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2944
timestamp 1018054153
transform 1 0 2352 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2946
timestamp 1018054153
transform 1 0 2368 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2948
timestamp 1018054153
transform 1 0 2384 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2950
timestamp 1018054153
transform 1 0 2400 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2952
timestamp 1018054153
transform 1 0 2416 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2954
timestamp 1018054153
transform 1 0 2432 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2956
timestamp 1018054153
transform 1 0 2448 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2958
timestamp 1018054153
transform 1 0 2464 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2960
timestamp 1018054153
transform 1 0 2480 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2962
timestamp 1018054153
transform 1 0 2496 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2964
timestamp 1018054153
transform 1 0 2512 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2966
timestamp 1018054153
transform 1 0 2528 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2968
timestamp 1018054153
transform 1 0 2544 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2970
timestamp 1018054153
transform 1 0 2560 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2972
timestamp 1018054153
transform 1 0 2576 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2974
timestamp 1018054153
transform 1 0 2592 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2976
timestamp 1018054153
transform 1 0 2608 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2978
timestamp 1018054153
transform 1 0 2624 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2980
timestamp 1018054153
transform 1 0 2640 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2982
timestamp 1018054153
transform 1 0 2656 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2984
timestamp 1018054153
transform 1 0 2672 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2986
timestamp 1018054153
transform 1 0 2688 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2988
timestamp 1018054153
transform 1 0 2704 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2990
timestamp 1018054153
transform 1 0 2720 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2992
timestamp 1018054153
transform 1 0 2736 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2994
timestamp 1018054153
transform 1 0 2752 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2996
timestamp 1018054153
transform 1 0 2768 0 -1 5680
box -16 -6 32 210
use FILL  FILL_2998
timestamp 1018054153
transform 1 0 2784 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3000
timestamp 1018054153
transform 1 0 2800 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3002
timestamp 1018054153
transform 1 0 2816 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3004
timestamp 1018054153
transform 1 0 2832 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3006
timestamp 1018054153
transform 1 0 2848 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3008
timestamp 1018054153
transform 1 0 2864 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3010
timestamp 1018054153
transform 1 0 2880 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3012
timestamp 1018054153
transform 1 0 2896 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3014
timestamp 1018054153
transform 1 0 2912 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3016
timestamp 1018054153
transform 1 0 2928 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3018
timestamp 1018054153
transform 1 0 2944 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3020
timestamp 1018054153
transform 1 0 2960 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3022
timestamp 1018054153
transform 1 0 2976 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3024
timestamp 1018054153
transform 1 0 2992 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3026
timestamp 1018054153
transform 1 0 3008 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3028
timestamp 1018054153
transform 1 0 3024 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3030
timestamp 1018054153
transform 1 0 3040 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3032
timestamp 1018054153
transform 1 0 3056 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3034
timestamp 1018054153
transform 1 0 3072 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3036
timestamp 1018054153
transform 1 0 3088 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3038
timestamp 1018054153
transform 1 0 3104 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3040
timestamp 1018054153
transform 1 0 3120 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3042
timestamp 1018054153
transform 1 0 3136 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3044
timestamp 1018054153
transform 1 0 3152 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3046
timestamp 1018054153
transform 1 0 3168 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3048
timestamp 1018054153
transform 1 0 3184 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3050
timestamp 1018054153
transform 1 0 3200 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3052
timestamp 1018054153
transform 1 0 3216 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3054
timestamp 1018054153
transform 1 0 3232 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3056
timestamp 1018054153
transform 1 0 3248 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3058
timestamp 1018054153
transform 1 0 3264 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3060
timestamp 1018054153
transform 1 0 3280 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3062
timestamp 1018054153
transform 1 0 3296 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3064
timestamp 1018054153
transform 1 0 3312 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3066
timestamp 1018054153
transform 1 0 3328 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3068
timestamp 1018054153
transform 1 0 3344 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3070
timestamp 1018054153
transform 1 0 3360 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3072
timestamp 1018054153
transform 1 0 3376 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3074
timestamp 1018054153
transform 1 0 3392 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3076
timestamp 1018054153
transform 1 0 3408 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3078
timestamp 1018054153
transform 1 0 3424 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3080
timestamp 1018054153
transform 1 0 3440 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3082
timestamp 1018054153
transform 1 0 3456 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3084
timestamp 1018054153
transform 1 0 3472 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3086
timestamp 1018054153
transform 1 0 3488 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3088
timestamp 1018054153
transform 1 0 3504 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3089
timestamp 1018054153
transform 1 0 3520 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3090
timestamp 1018054153
transform 1 0 3536 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3091
timestamp 1018054153
transform 1 0 3552 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3093
timestamp 1018054153
transform 1 0 3568 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3095
timestamp 1018054153
transform 1 0 3584 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3097
timestamp 1018054153
transform 1 0 3600 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3099
timestamp 1018054153
transform 1 0 3616 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3101
timestamp 1018054153
transform 1 0 3632 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3103
timestamp 1018054153
transform 1 0 3648 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3105
timestamp 1018054153
transform 1 0 3664 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3107
timestamp 1018054153
transform 1 0 3680 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3109
timestamp 1018054153
transform 1 0 3696 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3111
timestamp 1018054153
transform 1 0 3712 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3113
timestamp 1018054153
transform 1 0 3728 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3115
timestamp 1018054153
transform 1 0 3744 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3117
timestamp 1018054153
transform 1 0 3760 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3119
timestamp 1018054153
transform 1 0 3776 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3121
timestamp 1018054153
transform 1 0 3792 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3123
timestamp 1018054153
transform 1 0 3808 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3125
timestamp 1018054153
transform 1 0 3824 0 -1 5680
box -16 -6 32 210
use OAI21X1  OAI21X1_9
timestamp 1053722159
transform 1 0 3840 0 -1 5680
box -16 -6 68 210
use FILL  FILL_3131
timestamp 1018054153
transform 1 0 3904 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3133
timestamp 1018054153
transform 1 0 3920 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3135
timestamp 1018054153
transform 1 0 3936 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3137
timestamp 1018054153
transform 1 0 3952 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3139
timestamp 1018054153
transform 1 0 3968 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3141
timestamp 1018054153
transform 1 0 3984 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3143
timestamp 1018054153
transform 1 0 4000 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3145
timestamp 1018054153
transform 1 0 4016 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3147
timestamp 1018054153
transform 1 0 4032 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3149
timestamp 1018054153
transform 1 0 4048 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3151
timestamp 1018054153
transform 1 0 4064 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3153
timestamp 1018054153
transform 1 0 4080 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3155
timestamp 1018054153
transform 1 0 4096 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3157
timestamp 1018054153
transform 1 0 4112 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3159
timestamp 1018054153
transform 1 0 4128 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3161
timestamp 1018054153
transform 1 0 4144 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3163
timestamp 1018054153
transform 1 0 4160 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3165
timestamp 1018054153
transform 1 0 4176 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3167
timestamp 1018054153
transform 1 0 4192 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3169
timestamp 1018054153
transform 1 0 4208 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3171
timestamp 1018054153
transform 1 0 4224 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3173
timestamp 1018054153
transform 1 0 4240 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3175
timestamp 1018054153
transform 1 0 4256 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3177
timestamp 1018054153
transform 1 0 4272 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3179
timestamp 1018054153
transform 1 0 4288 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3181
timestamp 1018054153
transform 1 0 4304 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3183
timestamp 1018054153
transform 1 0 4320 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3185
timestamp 1018054153
transform 1 0 4336 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3187
timestamp 1018054153
transform 1 0 4352 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3189
timestamp 1018054153
transform 1 0 4368 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3191
timestamp 1018054153
transform 1 0 4384 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3193
timestamp 1018054153
transform 1 0 4400 0 -1 5680
box -16 -6 32 210
use AOI22X1  AOI22X1_0
timestamp 1053022145
transform 1 0 4416 0 -1 5680
box -16 -6 92 210
use FILL  FILL_3196
timestamp 1018054153
transform 1 0 4496 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3198
timestamp 1018054153
transform 1 0 4512 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3200
timestamp 1018054153
transform 1 0 4528 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3202
timestamp 1018054153
transform 1 0 4544 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3204
timestamp 1018054153
transform 1 0 4560 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3206
timestamp 1018054153
transform 1 0 4576 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3208
timestamp 1018054153
transform 1 0 4592 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3210
timestamp 1018054153
transform 1 0 4608 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3212
timestamp 1018054153
transform 1 0 4624 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3214
timestamp 1018054153
transform 1 0 4640 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3216
timestamp 1018054153
transform 1 0 4656 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3218
timestamp 1018054153
transform 1 0 4672 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3220
timestamp 1018054153
transform 1 0 4688 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3222
timestamp 1018054153
transform 1 0 4704 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3224
timestamp 1018054153
transform 1 0 4720 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3226
timestamp 1018054153
transform 1 0 4736 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3228
timestamp 1018054153
transform 1 0 4752 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3230
timestamp 1018054153
transform 1 0 4768 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3231
timestamp 1018054153
transform 1 0 4784 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3232
timestamp 1018054153
transform 1 0 4800 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3233
timestamp 1018054153
transform 1 0 4816 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3235
timestamp 1018054153
transform 1 0 4832 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3237
timestamp 1018054153
transform 1 0 4848 0 -1 5680
box -16 -6 32 210
use M3_M2  M3_M2_54
timestamp 1542725905
transform 1 0 4888 0 1 5490
box -6 -6 6 6
use FILL  FILL_3239
timestamp 1018054153
transform 1 0 4864 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3241
timestamp 1018054153
transform 1 0 4880 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3246
timestamp 1018054153
transform 1 0 4896 0 -1 5680
box -16 -6 32 210
use INVX1  INVX1_6
timestamp 1053022145
transform -1 0 4944 0 -1 5680
box -18 -6 52 210
use FILL  FILL_3247
timestamp 1018054153
transform 1 0 4944 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3249
timestamp 1018054153
transform 1 0 4960 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3251
timestamp 1018054153
transform 1 0 4976 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3253
timestamp 1018054153
transform 1 0 4992 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3255
timestamp 1018054153
transform 1 0 5008 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3257
timestamp 1018054153
transform 1 0 5024 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3260
timestamp 1018054153
transform 1 0 5040 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3261
timestamp 1018054153
transform 1 0 5056 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3262
timestamp 1018054153
transform 1 0 5072 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3263
timestamp 1018054153
transform 1 0 5088 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3264
timestamp 1018054153
transform 1 0 5104 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3265
timestamp 1018054153
transform 1 0 5120 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3266
timestamp 1018054153
transform 1 0 5136 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3267
timestamp 1018054153
transform 1 0 5152 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3268
timestamp 1018054153
transform 1 0 5168 0 -1 5680
box -16 -6 32 210
use NAND2X1  NAND2X1_8
timestamp 1053022145
transform 1 0 5184 0 -1 5680
box -16 -6 64 210
use FILL  FILL_3273
timestamp 1018054153
transform 1 0 5232 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3275
timestamp 1018054153
transform 1 0 5248 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3277
timestamp 1018054153
transform 1 0 5264 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3279
timestamp 1018054153
transform 1 0 5280 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3281
timestamp 1018054153
transform 1 0 5296 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3283
timestamp 1018054153
transform 1 0 5312 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3285
timestamp 1018054153
transform 1 0 5328 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3287
timestamp 1018054153
transform 1 0 5344 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3289
timestamp 1018054153
transform 1 0 5360 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3291
timestamp 1018054153
transform 1 0 5376 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3292
timestamp 1018054153
transform 1 0 5392 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3293
timestamp 1018054153
transform 1 0 5408 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3294
timestamp 1018054153
transform 1 0 5424 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3295
timestamp 1018054153
transform 1 0 5440 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3296
timestamp 1018054153
transform 1 0 5456 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3297
timestamp 1018054153
transform 1 0 5472 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3298
timestamp 1018054153
transform 1 0 5488 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3299
timestamp 1018054153
transform 1 0 5504 0 -1 5680
box -16 -6 32 210
use NAND2X1  NAND2X1_9
timestamp 1053022145
transform -1 0 5568 0 -1 5680
box -16 -6 64 210
use FILL  FILL_3300
timestamp 1018054153
transform 1 0 5568 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3301
timestamp 1018054153
transform 1 0 5584 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3302
timestamp 1018054153
transform 1 0 5600 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3303
timestamp 1018054153
transform 1 0 5616 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3305
timestamp 1018054153
transform 1 0 5632 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3307
timestamp 1018054153
transform 1 0 5648 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3309
timestamp 1018054153
transform 1 0 5664 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3311
timestamp 1018054153
transform 1 0 5680 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3313
timestamp 1018054153
transform 1 0 5696 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3315
timestamp 1018054153
transform 1 0 5712 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3317
timestamp 1018054153
transform 1 0 5728 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3319
timestamp 1018054153
transform 1 0 5744 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3321
timestamp 1018054153
transform 1 0 5760 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3323
timestamp 1018054153
transform 1 0 5776 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3325
timestamp 1018054153
transform 1 0 5792 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3327
timestamp 1018054153
transform 1 0 5808 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3329
timestamp 1018054153
transform 1 0 5824 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3331
timestamp 1018054153
transform 1 0 5840 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3337
timestamp 1018054153
transform 1 0 5856 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3338
timestamp 1018054153
transform 1 0 5872 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3339
timestamp 1018054153
transform 1 0 5888 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3340
timestamp 1018054153
transform 1 0 5904 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3341
timestamp 1018054153
transform 1 0 5920 0 -1 5680
box -16 -6 32 210
use NOR2X1  NOR2X1_6
timestamp 1053022145
transform -1 0 5984 0 -1 5680
box -16 -6 64 210
use FILL  FILL_3342
timestamp 1018054153
transform 1 0 5984 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3344
timestamp 1018054153
transform 1 0 6000 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3346
timestamp 1018054153
transform 1 0 6016 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3348
timestamp 1018054153
transform 1 0 6032 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3350
timestamp 1018054153
transform 1 0 6048 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3352
timestamp 1018054153
transform 1 0 6064 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3354
timestamp 1018054153
transform 1 0 6080 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3356
timestamp 1018054153
transform 1 0 6096 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3358
timestamp 1018054153
transform 1 0 6112 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3360
timestamp 1018054153
transform 1 0 6128 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3362
timestamp 1018054153
transform 1 0 6144 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3364
timestamp 1018054153
transform 1 0 6160 0 -1 5680
box -16 -6 32 210
use INVX1  INVX1_8
timestamp 1053022145
transform 1 0 6176 0 -1 5680
box -18 -6 52 210
use FILL  FILL_3367
timestamp 1018054153
transform 1 0 6208 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3368
timestamp 1018054153
transform 1 0 6224 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3370
timestamp 1018054153
transform 1 0 6240 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3372
timestamp 1018054153
transform 1 0 6256 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3374
timestamp 1018054153
transform 1 0 6272 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3376
timestamp 1018054153
transform 1 0 6288 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3378
timestamp 1018054153
transform 1 0 6304 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3380
timestamp 1018054153
transform 1 0 6320 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3382
timestamp 1018054153
transform 1 0 6336 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3384
timestamp 1018054153
transform 1 0 6352 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3386
timestamp 1018054153
transform 1 0 6368 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3388
timestamp 1018054153
transform 1 0 6384 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3390
timestamp 1018054153
transform 1 0 6400 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3392
timestamp 1018054153
transform 1 0 6416 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3394
timestamp 1018054153
transform 1 0 6432 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3396
timestamp 1018054153
transform 1 0 6448 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3401
timestamp 1018054153
transform 1 0 6464 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3402
timestamp 1018054153
transform 1 0 6480 0 -1 5680
box -16 -6 32 210
use AOI21X1  AOI21X1_2
timestamp 1090541997
transform 1 0 6496 0 -1 5680
box -14 -6 78 210
use FILL  FILL_3403
timestamp 1018054153
transform 1 0 6560 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3405
timestamp 1018054153
transform 1 0 6576 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3407
timestamp 1018054153
transform 1 0 6592 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3409
timestamp 1018054153
transform 1 0 6608 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3411
timestamp 1018054153
transform 1 0 6624 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3413
timestamp 1018054153
transform 1 0 6640 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3415
timestamp 1018054153
transform 1 0 6656 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3417
timestamp 1018054153
transform 1 0 6672 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3419
timestamp 1018054153
transform 1 0 6688 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3421
timestamp 1018054153
transform 1 0 6704 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3423
timestamp 1018054153
transform 1 0 6720 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3425
timestamp 1018054153
transform 1 0 6736 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3427
timestamp 1018054153
transform 1 0 6752 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3429
timestamp 1018054153
transform 1 0 6768 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3431
timestamp 1018054153
transform 1 0 6784 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3433
timestamp 1018054153
transform 1 0 6800 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3435
timestamp 1018054153
transform 1 0 6816 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3437
timestamp 1018054153
transform 1 0 6832 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3439
timestamp 1018054153
transform 1 0 6848 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3441
timestamp 1018054153
transform 1 0 6864 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3443
timestamp 1018054153
transform 1 0 6880 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3445
timestamp 1018054153
transform 1 0 6896 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3447
timestamp 1018054153
transform 1 0 6912 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3449
timestamp 1018054153
transform 1 0 6928 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3451
timestamp 1018054153
transform 1 0 6944 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3453
timestamp 1018054153
transform 1 0 6960 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3455
timestamp 1018054153
transform 1 0 6976 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3457
timestamp 1018054153
transform 1 0 6992 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3459
timestamp 1018054153
transform 1 0 7008 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3461
timestamp 1018054153
transform 1 0 7024 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3463
timestamp 1018054153
transform 1 0 7040 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3465
timestamp 1018054153
transform 1 0 7056 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3467
timestamp 1018054153
transform 1 0 7072 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3469
timestamp 1018054153
transform 1 0 7088 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3471
timestamp 1018054153
transform 1 0 7104 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3473
timestamp 1018054153
transform 1 0 7120 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3475
timestamp 1018054153
transform 1 0 7136 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3477
timestamp 1018054153
transform 1 0 7152 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3479
timestamp 1018054153
transform 1 0 7168 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3481
timestamp 1018054153
transform 1 0 7184 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3483
timestamp 1018054153
transform 1 0 7200 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3485
timestamp 1018054153
transform 1 0 7216 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3487
timestamp 1018054153
transform 1 0 7232 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3489
timestamp 1018054153
transform 1 0 7248 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3491
timestamp 1018054153
transform 1 0 7264 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3493
timestamp 1018054153
transform 1 0 7280 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3495
timestamp 1018054153
transform 1 0 7296 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3497
timestamp 1018054153
transform 1 0 7312 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3499
timestamp 1018054153
transform 1 0 7328 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3501
timestamp 1018054153
transform 1 0 7344 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3503
timestamp 1018054153
transform 1 0 7360 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3505
timestamp 1018054153
transform 1 0 7376 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3507
timestamp 1018054153
transform 1 0 7392 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3509
timestamp 1018054153
transform 1 0 7408 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3511
timestamp 1018054153
transform 1 0 7424 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3513
timestamp 1018054153
transform 1 0 7440 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3515
timestamp 1018054153
transform 1 0 7456 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3517
timestamp 1018054153
transform 1 0 7472 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3519
timestamp 1018054153
transform 1 0 7488 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3521
timestamp 1018054153
transform 1 0 7504 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3523
timestamp 1018054153
transform 1 0 7520 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3525
timestamp 1018054153
transform 1 0 7536 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3527
timestamp 1018054153
transform 1 0 7552 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3529
timestamp 1018054153
transform 1 0 7568 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3531
timestamp 1018054153
transform 1 0 7584 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3533
timestamp 1018054153
transform 1 0 7600 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3535
timestamp 1018054153
transform 1 0 7616 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3537
timestamp 1018054153
transform 1 0 7632 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3539
timestamp 1018054153
transform 1 0 7648 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3541
timestamp 1018054153
transform 1 0 7664 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3543
timestamp 1018054153
transform 1 0 7680 0 -1 5680
box -16 -6 32 210
use FILL  FILL_3545
timestamp 1018054153
transform 1 0 7696 0 -1 5680
box -16 -6 32 210
use PADNC  PADNC_7
timestamp 1084294400
transform 0 1 8000 -1 0 6200
box -6 -6 606 2000
use M3_M2  M3_M2_53
timestamp 1542725905
transform 1 0 8002 0 1 5510
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_19
timestamp 1542725905
transform 1 0 7788 0 1 5480
box -48 -6 48 6
use FILL  FILL_3547
timestamp 1018054153
transform 1 0 7712 0 -1 5680
box -16 -6 32 210
use M2_M1  M2_M1_165
timestamp 1542725905
transform 1 0 4056 0 1 5350
box -4 -4 4 4
use M3_M2  M3_M2_55
timestamp 1542725905
transform 1 0 4184 0 1 5450
box -6 -6 6 6
use M2_M1  M2_M1_174
timestamp 1542725905
transform 1 0 4216 0 1 5330
box -4 -4 4 4
use M2_M1  M2_M1_166
timestamp 1542725905
transform 1 0 4408 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_175
timestamp 1542725905
transform 1 0 4488 0 1 5330
box -4 -4 4 4
use M3_M2  M3_M2_56
timestamp 1542725905
transform 1 0 4536 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_157
timestamp 1542725905
transform 1 0 4536 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_158
timestamp 1542725905
transform 1 0 4552 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_176
timestamp 1542725905
transform 1 0 4792 0 1 5330
box -4 -4 4 4
use M2_M1  M2_M1_167
timestamp 1542725905
transform 1 0 4968 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_159
timestamp 1542725905
transform 1 0 5048 0 1 5370
box -4 -4 4 4
use M3_M2  M3_M2_57
timestamp 1542725905
transform 1 0 5160 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_160
timestamp 1542725905
transform 1 0 5144 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_168
timestamp 1542725905
transform 1 0 5160 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_177
timestamp 1542725905
transform 1 0 5256 0 1 5330
box -4 -4 4 4
use M3_M2  M3_M2_58
timestamp 1542725905
transform 1 0 5336 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_169
timestamp 1542725905
transform 1 0 5512 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_178
timestamp 1542725905
transform 1 0 5496 0 1 5330
box -4 -4 4 4
use M3_M2  M3_M2_59
timestamp 1542725905
transform 1 0 5560 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_161
timestamp 1542725905
transform 1 0 5544 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_179
timestamp 1542725905
transform 1 0 5720 0 1 5330
box -4 -4 4 4
use M2_M1  M2_M1_170
timestamp 1542725905
transform 1 0 5752 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_180
timestamp 1542725905
transform 1 0 5784 0 1 5330
box -4 -4 4 4
use M2_M1  M2_M1_171
timestamp 1542725905
transform 1 0 5864 0 1 5350
box -4 -4 4 4
use M3_M2  M3_M2_60
timestamp 1542725905
transform 1 0 6152 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_172
timestamp 1542725905
transform 1 0 6264 0 1 5350
box -4 -4 4 4
use M3_M2  M3_M2_62
timestamp 1542725905
transform 1 0 6264 0 1 5330
box -6 -6 6 6
use M3_M2  M3_M2_61
timestamp 1542725905
transform 1 0 6328 0 1 5390
box -6 -6 6 6
use M2_M1  M2_M1_162
timestamp 1542725905
transform 1 0 6328 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_173
timestamp 1542725905
transform 1 0 6600 0 1 5350
box -4 -4 4 4
use M2_M1  M2_M1_163
timestamp 1542725905
transform 1 0 6792 0 1 5370
box -4 -4 4 4
use M2_M1  M2_M1_164
timestamp 1542725905
transform 1 0 6824 0 1 5370
box -4 -4 4 4
use M3_M2  M3_M2_63
timestamp 1542725905
transform 1 0 6792 0 1 5330
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_20
timestamp 1542725905
transform 1 0 2092 0 1 5280
box -48 -6 48 6
use FILL  FILL_3548
timestamp 1018054153
transform 1 0 2272 0 1 5280
box -16 -6 32 210
use FILL  FILL_3550
timestamp 1018054153
transform 1 0 2288 0 1 5280
box -16 -6 32 210
use FILL  FILL_3552
timestamp 1018054153
transform 1 0 2304 0 1 5280
box -16 -6 32 210
use FILL  FILL_3554
timestamp 1018054153
transform 1 0 2320 0 1 5280
box -16 -6 32 210
use FILL  FILL_3556
timestamp 1018054153
transform 1 0 2336 0 1 5280
box -16 -6 32 210
use FILL  FILL_3558
timestamp 1018054153
transform 1 0 2352 0 1 5280
box -16 -6 32 210
use FILL  FILL_3560
timestamp 1018054153
transform 1 0 2368 0 1 5280
box -16 -6 32 210
use FILL  FILL_3562
timestamp 1018054153
transform 1 0 2384 0 1 5280
box -16 -6 32 210
use FILL  FILL_3564
timestamp 1018054153
transform 1 0 2400 0 1 5280
box -16 -6 32 210
use FILL  FILL_3566
timestamp 1018054153
transform 1 0 2416 0 1 5280
box -16 -6 32 210
use FILL  FILL_3568
timestamp 1018054153
transform 1 0 2432 0 1 5280
box -16 -6 32 210
use FILL  FILL_3570
timestamp 1018054153
transform 1 0 2448 0 1 5280
box -16 -6 32 210
use FILL  FILL_3572
timestamp 1018054153
transform 1 0 2464 0 1 5280
box -16 -6 32 210
use FILL  FILL_3574
timestamp 1018054153
transform 1 0 2480 0 1 5280
box -16 -6 32 210
use FILL  FILL_3576
timestamp 1018054153
transform 1 0 2496 0 1 5280
box -16 -6 32 210
use FILL  FILL_3578
timestamp 1018054153
transform 1 0 2512 0 1 5280
box -16 -6 32 210
use FILL  FILL_3580
timestamp 1018054153
transform 1 0 2528 0 1 5280
box -16 -6 32 210
use FILL  FILL_3582
timestamp 1018054153
transform 1 0 2544 0 1 5280
box -16 -6 32 210
use FILL  FILL_3584
timestamp 1018054153
transform 1 0 2560 0 1 5280
box -16 -6 32 210
use FILL  FILL_3586
timestamp 1018054153
transform 1 0 2576 0 1 5280
box -16 -6 32 210
use FILL  FILL_3588
timestamp 1018054153
transform 1 0 2592 0 1 5280
box -16 -6 32 210
use FILL  FILL_3590
timestamp 1018054153
transform 1 0 2608 0 1 5280
box -16 -6 32 210
use FILL  FILL_3592
timestamp 1018054153
transform 1 0 2624 0 1 5280
box -16 -6 32 210
use FILL  FILL_3594
timestamp 1018054153
transform 1 0 2640 0 1 5280
box -16 -6 32 210
use FILL  FILL_3596
timestamp 1018054153
transform 1 0 2656 0 1 5280
box -16 -6 32 210
use FILL  FILL_3598
timestamp 1018054153
transform 1 0 2672 0 1 5280
box -16 -6 32 210
use FILL  FILL_3600
timestamp 1018054153
transform 1 0 2688 0 1 5280
box -16 -6 32 210
use FILL  FILL_3602
timestamp 1018054153
transform 1 0 2704 0 1 5280
box -16 -6 32 210
use FILL  FILL_3604
timestamp 1018054153
transform 1 0 2720 0 1 5280
box -16 -6 32 210
use FILL  FILL_3606
timestamp 1018054153
transform 1 0 2736 0 1 5280
box -16 -6 32 210
use FILL  FILL_3608
timestamp 1018054153
transform 1 0 2752 0 1 5280
box -16 -6 32 210
use FILL  FILL_3610
timestamp 1018054153
transform 1 0 2768 0 1 5280
box -16 -6 32 210
use FILL  FILL_3612
timestamp 1018054153
transform 1 0 2784 0 1 5280
box -16 -6 32 210
use FILL  FILL_3614
timestamp 1018054153
transform 1 0 2800 0 1 5280
box -16 -6 32 210
use FILL  FILL_3616
timestamp 1018054153
transform 1 0 2816 0 1 5280
box -16 -6 32 210
use FILL  FILL_3618
timestamp 1018054153
transform 1 0 2832 0 1 5280
box -16 -6 32 210
use FILL  FILL_3620
timestamp 1018054153
transform 1 0 2848 0 1 5280
box -16 -6 32 210
use FILL  FILL_3622
timestamp 1018054153
transform 1 0 2864 0 1 5280
box -16 -6 32 210
use FILL  FILL_3624
timestamp 1018054153
transform 1 0 2880 0 1 5280
box -16 -6 32 210
use FILL  FILL_3626
timestamp 1018054153
transform 1 0 2896 0 1 5280
box -16 -6 32 210
use FILL  FILL_3628
timestamp 1018054153
transform 1 0 2912 0 1 5280
box -16 -6 32 210
use FILL  FILL_3630
timestamp 1018054153
transform 1 0 2928 0 1 5280
box -16 -6 32 210
use FILL  FILL_3632
timestamp 1018054153
transform 1 0 2944 0 1 5280
box -16 -6 32 210
use FILL  FILL_3634
timestamp 1018054153
transform 1 0 2960 0 1 5280
box -16 -6 32 210
use FILL  FILL_3636
timestamp 1018054153
transform 1 0 2976 0 1 5280
box -16 -6 32 210
use FILL  FILL_3638
timestamp 1018054153
transform 1 0 2992 0 1 5280
box -16 -6 32 210
use FILL  FILL_3640
timestamp 1018054153
transform 1 0 3008 0 1 5280
box -16 -6 32 210
use FILL  FILL_3642
timestamp 1018054153
transform 1 0 3024 0 1 5280
box -16 -6 32 210
use FILL  FILL_3644
timestamp 1018054153
transform 1 0 3040 0 1 5280
box -16 -6 32 210
use FILL  FILL_3646
timestamp 1018054153
transform 1 0 3056 0 1 5280
box -16 -6 32 210
use FILL  FILL_3648
timestamp 1018054153
transform 1 0 3072 0 1 5280
box -16 -6 32 210
use FILL  FILL_3650
timestamp 1018054153
transform 1 0 3088 0 1 5280
box -16 -6 32 210
use FILL  FILL_3652
timestamp 1018054153
transform 1 0 3104 0 1 5280
box -16 -6 32 210
use FILL  FILL_3654
timestamp 1018054153
transform 1 0 3120 0 1 5280
box -16 -6 32 210
use FILL  FILL_3656
timestamp 1018054153
transform 1 0 3136 0 1 5280
box -16 -6 32 210
use FILL  FILL_3658
timestamp 1018054153
transform 1 0 3152 0 1 5280
box -16 -6 32 210
use FILL  FILL_3660
timestamp 1018054153
transform 1 0 3168 0 1 5280
box -16 -6 32 210
use FILL  FILL_3662
timestamp 1018054153
transform 1 0 3184 0 1 5280
box -16 -6 32 210
use FILL  FILL_3664
timestamp 1018054153
transform 1 0 3200 0 1 5280
box -16 -6 32 210
use FILL  FILL_3666
timestamp 1018054153
transform 1 0 3216 0 1 5280
box -16 -6 32 210
use FILL  FILL_3668
timestamp 1018054153
transform 1 0 3232 0 1 5280
box -16 -6 32 210
use FILL  FILL_3670
timestamp 1018054153
transform 1 0 3248 0 1 5280
box -16 -6 32 210
use FILL  FILL_3672
timestamp 1018054153
transform 1 0 3264 0 1 5280
box -16 -6 32 210
use FILL  FILL_3674
timestamp 1018054153
transform 1 0 3280 0 1 5280
box -16 -6 32 210
use FILL  FILL_3676
timestamp 1018054153
transform 1 0 3296 0 1 5280
box -16 -6 32 210
use FILL  FILL_3678
timestamp 1018054153
transform 1 0 3312 0 1 5280
box -16 -6 32 210
use FILL  FILL_3680
timestamp 1018054153
transform 1 0 3328 0 1 5280
box -16 -6 32 210
use FILL  FILL_3682
timestamp 1018054153
transform 1 0 3344 0 1 5280
box -16 -6 32 210
use FILL  FILL_3684
timestamp 1018054153
transform 1 0 3360 0 1 5280
box -16 -6 32 210
use FILL  FILL_3686
timestamp 1018054153
transform 1 0 3376 0 1 5280
box -16 -6 32 210
use FILL  FILL_3688
timestamp 1018054153
transform 1 0 3392 0 1 5280
box -16 -6 32 210
use FILL  FILL_3690
timestamp 1018054153
transform 1 0 3408 0 1 5280
box -16 -6 32 210
use FILL  FILL_3692
timestamp 1018054153
transform 1 0 3424 0 1 5280
box -16 -6 32 210
use FILL  FILL_3694
timestamp 1018054153
transform 1 0 3440 0 1 5280
box -16 -6 32 210
use FILL  FILL_3696
timestamp 1018054153
transform 1 0 3456 0 1 5280
box -16 -6 32 210
use FILL  FILL_3698
timestamp 1018054153
transform 1 0 3472 0 1 5280
box -16 -6 32 210
use FILL  FILL_3700
timestamp 1018054153
transform 1 0 3488 0 1 5280
box -16 -6 32 210
use FILL  FILL_3702
timestamp 1018054153
transform 1 0 3504 0 1 5280
box -16 -6 32 210
use FILL  FILL_3704
timestamp 1018054153
transform 1 0 3520 0 1 5280
box -16 -6 32 210
use FILL  FILL_3706
timestamp 1018054153
transform 1 0 3536 0 1 5280
box -16 -6 32 210
use FILL  FILL_3708
timestamp 1018054153
transform 1 0 3552 0 1 5280
box -16 -6 32 210
use FILL  FILL_3710
timestamp 1018054153
transform 1 0 3568 0 1 5280
box -16 -6 32 210
use FILL  FILL_3712
timestamp 1018054153
transform 1 0 3584 0 1 5280
box -16 -6 32 210
use FILL  FILL_3714
timestamp 1018054153
transform 1 0 3600 0 1 5280
box -16 -6 32 210
use FILL  FILL_3716
timestamp 1018054153
transform 1 0 3616 0 1 5280
box -16 -6 32 210
use FILL  FILL_3718
timestamp 1018054153
transform 1 0 3632 0 1 5280
box -16 -6 32 210
use FILL  FILL_3720
timestamp 1018054153
transform 1 0 3648 0 1 5280
box -16 -6 32 210
use FILL  FILL_3722
timestamp 1018054153
transform 1 0 3664 0 1 5280
box -16 -6 32 210
use FILL  FILL_3724
timestamp 1018054153
transform 1 0 3680 0 1 5280
box -16 -6 32 210
use FILL  FILL_3726
timestamp 1018054153
transform 1 0 3696 0 1 5280
box -16 -6 32 210
use FILL  FILL_3728
timestamp 1018054153
transform 1 0 3712 0 1 5280
box -16 -6 32 210
use FILL  FILL_3730
timestamp 1018054153
transform 1 0 3728 0 1 5280
box -16 -6 32 210
use FILL  FILL_3732
timestamp 1018054153
transform 1 0 3744 0 1 5280
box -16 -6 32 210
use FILL  FILL_3734
timestamp 1018054153
transform 1 0 3760 0 1 5280
box -16 -6 32 210
use FILL  FILL_3736
timestamp 1018054153
transform 1 0 3776 0 1 5280
box -16 -6 32 210
use FILL  FILL_3738
timestamp 1018054153
transform 1 0 3792 0 1 5280
box -16 -6 32 210
use FILL  FILL_3740
timestamp 1018054153
transform 1 0 3808 0 1 5280
box -16 -6 32 210
use FILL  FILL_3742
timestamp 1018054153
transform 1 0 3824 0 1 5280
box -16 -6 32 210
use FILL  FILL_3744
timestamp 1018054153
transform 1 0 3840 0 1 5280
box -16 -6 32 210
use FILL  FILL_3746
timestamp 1018054153
transform 1 0 3856 0 1 5280
box -16 -6 32 210
use FILL  FILL_3748
timestamp 1018054153
transform 1 0 3872 0 1 5280
box -16 -6 32 210
use FILL  FILL_3750
timestamp 1018054153
transform 1 0 3888 0 1 5280
box -16 -6 32 210
use FILL  FILL_3752
timestamp 1018054153
transform 1 0 3904 0 1 5280
box -16 -6 32 210
use FILL  FILL_3754
timestamp 1018054153
transform 1 0 3920 0 1 5280
box -16 -6 32 210
use FILL  FILL_3756
timestamp 1018054153
transform 1 0 3936 0 1 5280
box -16 -6 32 210
use FILL  FILL_3758
timestamp 1018054153
transform 1 0 3952 0 1 5280
box -16 -6 32 210
use FILL  FILL_3760
timestamp 1018054153
transform 1 0 3968 0 1 5280
box -16 -6 32 210
use FILL  FILL_3762
timestamp 1018054153
transform 1 0 3984 0 1 5280
box -16 -6 32 210
use FILL  FILL_3764
timestamp 1018054153
transform 1 0 4000 0 1 5280
box -16 -6 32 210
use FILL  FILL_3766
timestamp 1018054153
transform 1 0 4016 0 1 5280
box -16 -6 32 210
use FILL  FILL_3768
timestamp 1018054153
transform 1 0 4032 0 1 5280
box -16 -6 32 210
use FILL  FILL_3770
timestamp 1018054153
transform 1 0 4048 0 1 5280
box -16 -6 32 210
use FILL  FILL_3772
timestamp 1018054153
transform 1 0 4064 0 1 5280
box -16 -6 32 210
use FILL  FILL_3774
timestamp 1018054153
transform 1 0 4080 0 1 5280
box -16 -6 32 210
use FILL  FILL_3776
timestamp 1018054153
transform 1 0 4096 0 1 5280
box -16 -6 32 210
use FILL  FILL_3778
timestamp 1018054153
transform 1 0 4112 0 1 5280
box -16 -6 32 210
use FILL  FILL_3780
timestamp 1018054153
transform 1 0 4128 0 1 5280
box -16 -6 32 210
use FILL  FILL_3782
timestamp 1018054153
transform 1 0 4144 0 1 5280
box -16 -6 32 210
use FILL  FILL_3784
timestamp 1018054153
transform 1 0 4160 0 1 5280
box -16 -6 32 210
use FILL  FILL_3786
timestamp 1018054153
transform 1 0 4176 0 1 5280
box -16 -6 32 210
use FILL  FILL_3788
timestamp 1018054153
transform 1 0 4192 0 1 5280
box -16 -6 32 210
use INVX1  INVX1_9
timestamp 1053022145
transform 1 0 4208 0 1 5280
box -18 -6 52 210
use FILL  FILL_3790
timestamp 1018054153
transform 1 0 4240 0 1 5280
box -16 -6 32 210
use FILL  FILL_3794
timestamp 1018054153
transform 1 0 4256 0 1 5280
box -16 -6 32 210
use FILL  FILL_3796
timestamp 1018054153
transform 1 0 4272 0 1 5280
box -16 -6 32 210
use FILL  FILL_3798
timestamp 1018054153
transform 1 0 4288 0 1 5280
box -16 -6 32 210
use FILL  FILL_3800
timestamp 1018054153
transform 1 0 4304 0 1 5280
box -16 -6 32 210
use FILL  FILL_3802
timestamp 1018054153
transform 1 0 4320 0 1 5280
box -16 -6 32 210
use FILL  FILL_3804
timestamp 1018054153
transform 1 0 4336 0 1 5280
box -16 -6 32 210
use FILL  FILL_3806
timestamp 1018054153
transform 1 0 4352 0 1 5280
box -16 -6 32 210
use FILL  FILL_3808
timestamp 1018054153
transform 1 0 4368 0 1 5280
box -16 -6 32 210
use FILL  FILL_3810
timestamp 1018054153
transform 1 0 4384 0 1 5280
box -16 -6 32 210
use FILL  FILL_3811
timestamp 1018054153
transform 1 0 4400 0 1 5280
box -16 -6 32 210
use FILL  FILL_3812
timestamp 1018054153
transform 1 0 4416 0 1 5280
box -16 -6 32 210
use FILL  FILL_3814
timestamp 1018054153
transform 1 0 4432 0 1 5280
box -16 -6 32 210
use FILL  FILL_3816
timestamp 1018054153
transform 1 0 4448 0 1 5280
box -16 -6 32 210
use FILL  FILL_3818
timestamp 1018054153
transform 1 0 4464 0 1 5280
box -16 -6 32 210
use FILL  FILL_3820
timestamp 1018054153
transform 1 0 4480 0 1 5280
box -16 -6 32 210
use NOR2X1  NOR2X1_8
timestamp 1053022145
transform 1 0 4496 0 1 5280
box -16 -6 64 210
use FILL  FILL_3822
timestamp 1018054153
transform 1 0 4544 0 1 5280
box -16 -6 32 210
use FILL  FILL_3827
timestamp 1018054153
transform 1 0 4560 0 1 5280
box -16 -6 32 210
use FILL  FILL_3829
timestamp 1018054153
transform 1 0 4576 0 1 5280
box -16 -6 32 210
use FILL  FILL_3831
timestamp 1018054153
transform 1 0 4592 0 1 5280
box -16 -6 32 210
use FILL  FILL_3833
timestamp 1018054153
transform 1 0 4608 0 1 5280
box -16 -6 32 210
use FILL  FILL_3835
timestamp 1018054153
transform 1 0 4624 0 1 5280
box -16 -6 32 210
use FILL  FILL_3837
timestamp 1018054153
transform 1 0 4640 0 1 5280
box -16 -6 32 210
use FILL  FILL_3839
timestamp 1018054153
transform 1 0 4656 0 1 5280
box -16 -6 32 210
use FILL  FILL_3841
timestamp 1018054153
transform 1 0 4672 0 1 5280
box -16 -6 32 210
use FILL  FILL_3843
timestamp 1018054153
transform 1 0 4688 0 1 5280
box -16 -6 32 210
use FILL  FILL_3844
timestamp 1018054153
transform 1 0 4704 0 1 5280
box -16 -6 32 210
use FILL  FILL_3845
timestamp 1018054153
transform 1 0 4720 0 1 5280
box -16 -6 32 210
use FILL  FILL_3846
timestamp 1018054153
transform 1 0 4736 0 1 5280
box -16 -6 32 210
use NOR2X1  NOR2X1_9
timestamp 1053022145
transform -1 0 4800 0 1 5280
box -16 -6 64 210
use FILL  FILL_3847
timestamp 1018054153
transform 1 0 4800 0 1 5280
box -16 -6 32 210
use FILL  FILL_3852
timestamp 1018054153
transform 1 0 4816 0 1 5280
box -16 -6 32 210
use FILL  FILL_3854
timestamp 1018054153
transform 1 0 4832 0 1 5280
box -16 -6 32 210
use FILL  FILL_3856
timestamp 1018054153
transform 1 0 4848 0 1 5280
box -16 -6 32 210
use FILL  FILL_3858
timestamp 1018054153
transform 1 0 4864 0 1 5280
box -16 -6 32 210
use FILL  FILL_3860
timestamp 1018054153
transform 1 0 4880 0 1 5280
box -16 -6 32 210
use FILL  FILL_3862
timestamp 1018054153
transform 1 0 4896 0 1 5280
box -16 -6 32 210
use FILL  FILL_3864
timestamp 1018054153
transform 1 0 4912 0 1 5280
box -16 -6 32 210
use FILL  FILL_3866
timestamp 1018054153
transform 1 0 4928 0 1 5280
box -16 -6 32 210
use FILL  FILL_3868
timestamp 1018054153
transform 1 0 4944 0 1 5280
box -16 -6 32 210
use FILL  FILL_3870
timestamp 1018054153
transform 1 0 4960 0 1 5280
box -16 -6 32 210
use FILL  FILL_3872
timestamp 1018054153
transform 1 0 4976 0 1 5280
box -16 -6 32 210
use FILL  FILL_3873
timestamp 1018054153
transform 1 0 4992 0 1 5280
box -16 -6 32 210
use FILL  FILL_3874
timestamp 1018054153
transform 1 0 5008 0 1 5280
box -16 -6 32 210
use AND2X2  AND2X2_0
timestamp 1090541974
transform 1 0 5024 0 1 5280
box -16 -6 80 210
use FILL  FILL_3875
timestamp 1018054153
transform 1 0 5088 0 1 5280
box -16 -6 32 210
use FILL  FILL_3876
timestamp 1018054153
transform 1 0 5104 0 1 5280
box -16 -6 32 210
use FILL  FILL_3879
timestamp 1018054153
transform 1 0 5120 0 1 5280
box -16 -6 32 210
use FILL  FILL_3881
timestamp 1018054153
transform 1 0 5136 0 1 5280
box -16 -6 32 210
use FILL  FILL_3883
timestamp 1018054153
transform 1 0 5152 0 1 5280
box -16 -6 32 210
use FILL  FILL_3885
timestamp 1018054153
transform 1 0 5168 0 1 5280
box -16 -6 32 210
use FILL  FILL_3887
timestamp 1018054153
transform 1 0 5184 0 1 5280
box -16 -6 32 210
use FILL  FILL_3889
timestamp 1018054153
transform 1 0 5200 0 1 5280
box -16 -6 32 210
use FILL  FILL_3891
timestamp 1018054153
transform 1 0 5216 0 1 5280
box -16 -6 32 210
use FILL  FILL_3893
timestamp 1018054153
transform 1 0 5232 0 1 5280
box -16 -6 32 210
use FILL  FILL_3895
timestamp 1018054153
transform 1 0 5248 0 1 5280
box -16 -6 32 210
use FILL  FILL_3897
timestamp 1018054153
transform 1 0 5264 0 1 5280
box -16 -6 32 210
use INVX1  INVX1_11
timestamp 1053022145
transform 1 0 5280 0 1 5280
box -18 -6 52 210
use FILL  FILL_3899
timestamp 1018054153
transform 1 0 5312 0 1 5280
box -16 -6 32 210
use FILL  FILL_3903
timestamp 1018054153
transform 1 0 5328 0 1 5280
box -16 -6 32 210
use FILL  FILL_3904
timestamp 1018054153
transform 1 0 5344 0 1 5280
box -16 -6 32 210
use FILL  FILL_3905
timestamp 1018054153
transform 1 0 5360 0 1 5280
box -16 -6 32 210
use FILL  FILL_3907
timestamp 1018054153
transform 1 0 5376 0 1 5280
box -16 -6 32 210
use FILL  FILL_3909
timestamp 1018054153
transform 1 0 5392 0 1 5280
box -16 -6 32 210
use FILL  FILL_3911
timestamp 1018054153
transform 1 0 5408 0 1 5280
box -16 -6 32 210
use FILL  FILL_3913
timestamp 1018054153
transform 1 0 5424 0 1 5280
box -16 -6 32 210
use FILL  FILL_3915
timestamp 1018054153
transform 1 0 5440 0 1 5280
box -16 -6 32 210
use FILL  FILL_3917
timestamp 1018054153
transform 1 0 5456 0 1 5280
box -16 -6 32 210
use FILL  FILL_3919
timestamp 1018054153
transform 1 0 5472 0 1 5280
box -16 -6 32 210
use FILL  FILL_3921
timestamp 1018054153
transform 1 0 5488 0 1 5280
box -16 -6 32 210
use NOR2X1  NOR2X1_10
timestamp 1053022145
transform 1 0 5504 0 1 5280
box -16 -6 64 210
use FILL  FILL_3923
timestamp 1018054153
transform 1 0 5552 0 1 5280
box -16 -6 32 210
use FILL  FILL_3928
timestamp 1018054153
transform 1 0 5568 0 1 5280
box -16 -6 32 210
use FILL  FILL_3930
timestamp 1018054153
transform 1 0 5584 0 1 5280
box -16 -6 32 210
use FILL  FILL_3932
timestamp 1018054153
transform 1 0 5600 0 1 5280
box -16 -6 32 210
use FILL  FILL_3934
timestamp 1018054153
transform 1 0 5616 0 1 5280
box -16 -6 32 210
use FILL  FILL_3936
timestamp 1018054153
transform 1 0 5632 0 1 5280
box -16 -6 32 210
use FILL  FILL_3938
timestamp 1018054153
transform 1 0 5648 0 1 5280
box -16 -6 32 210
use FILL  FILL_3940
timestamp 1018054153
transform 1 0 5664 0 1 5280
box -16 -6 32 210
use FILL  FILL_3942
timestamp 1018054153
transform 1 0 5680 0 1 5280
box -16 -6 32 210
use FILL  FILL_3944
timestamp 1018054153
transform 1 0 5696 0 1 5280
box -16 -6 32 210
use FILL  FILL_3946
timestamp 1018054153
transform 1 0 5712 0 1 5280
box -16 -6 32 210
use FILL  FILL_3948
timestamp 1018054153
transform 1 0 5728 0 1 5280
box -16 -6 32 210
use INVX1  INVX1_13
timestamp 1053022145
transform 1 0 5744 0 1 5280
box -18 -6 52 210
use FILL  FILL_3950
timestamp 1018054153
transform 1 0 5776 0 1 5280
box -16 -6 32 210
use FILL  FILL_3954
timestamp 1018054153
transform 1 0 5792 0 1 5280
box -16 -6 32 210
use FILL  FILL_3956
timestamp 1018054153
transform 1 0 5808 0 1 5280
box -16 -6 32 210
use FILL  FILL_3958
timestamp 1018054153
transform 1 0 5824 0 1 5280
box -16 -6 32 210
use FILL  FILL_3960
timestamp 1018054153
transform 1 0 5840 0 1 5280
box -16 -6 32 210
use FILL  FILL_3962
timestamp 1018054153
transform 1 0 5856 0 1 5280
box -16 -6 32 210
use FILL  FILL_3964
timestamp 1018054153
transform 1 0 5872 0 1 5280
box -16 -6 32 210
use FILL  FILL_3966
timestamp 1018054153
transform 1 0 5888 0 1 5280
box -16 -6 32 210
use FILL  FILL_3968
timestamp 1018054153
transform 1 0 5904 0 1 5280
box -16 -6 32 210
use FILL  FILL_3970
timestamp 1018054153
transform 1 0 5920 0 1 5280
box -16 -6 32 210
use FILL  FILL_3971
timestamp 1018054153
transform 1 0 5936 0 1 5280
box -16 -6 32 210
use FILL  FILL_3972
timestamp 1018054153
transform 1 0 5952 0 1 5280
box -16 -6 32 210
use FILL  FILL_3973
timestamp 1018054153
transform 1 0 5968 0 1 5280
box -16 -6 32 210
use FILL  FILL_3974
timestamp 1018054153
transform 1 0 5984 0 1 5280
box -16 -6 32 210
use FILL  FILL_3975
timestamp 1018054153
transform 1 0 6000 0 1 5280
box -16 -6 32 210
use FILL  FILL_3976
timestamp 1018054153
transform 1 0 6016 0 1 5280
box -16 -6 32 210
use FILL  FILL_3977
timestamp 1018054153
transform 1 0 6032 0 1 5280
box -16 -6 32 210
use FILL  FILL_3979
timestamp 1018054153
transform 1 0 6048 0 1 5280
box -16 -6 32 210
use FILL  FILL_3981
timestamp 1018054153
transform 1 0 6064 0 1 5280
box -16 -6 32 210
use FILL  FILL_3983
timestamp 1018054153
transform 1 0 6080 0 1 5280
box -16 -6 32 210
use FILL  FILL_3985
timestamp 1018054153
transform 1 0 6096 0 1 5280
box -16 -6 32 210
use FILL  FILL_3987
timestamp 1018054153
transform 1 0 6112 0 1 5280
box -16 -6 32 210
use FILL  FILL_3989
timestamp 1018054153
transform 1 0 6128 0 1 5280
box -16 -6 32 210
use FILL  FILL_3991
timestamp 1018054153
transform 1 0 6144 0 1 5280
box -16 -6 32 210
use FILL  FILL_3993
timestamp 1018054153
transform 1 0 6160 0 1 5280
box -16 -6 32 210
use FILL  FILL_3995
timestamp 1018054153
transform 1 0 6176 0 1 5280
box -16 -6 32 210
use FILL  FILL_3997
timestamp 1018054153
transform 1 0 6192 0 1 5280
box -16 -6 32 210
use FILL  FILL_3999
timestamp 1018054153
transform 1 0 6208 0 1 5280
box -16 -6 32 210
use FILL  FILL_4001
timestamp 1018054153
transform 1 0 6224 0 1 5280
box -16 -6 32 210
use FILL  FILL_4003
timestamp 1018054153
transform 1 0 6240 0 1 5280
box -16 -6 32 210
use FILL  FILL_4005
timestamp 1018054153
transform 1 0 6256 0 1 5280
box -16 -6 32 210
use XOR2X1  XOR2X1_5
timestamp 1053359338
transform 1 0 6272 0 1 5280
box -16 -6 128 210
use FILL  FILL_4007
timestamp 1018054153
transform 1 0 6384 0 1 5280
box -16 -6 32 210
use FILL  FILL_4016
timestamp 1018054153
transform 1 0 6400 0 1 5280
box -16 -6 32 210
use FILL  FILL_4018
timestamp 1018054153
transform 1 0 6416 0 1 5280
box -16 -6 32 210
use FILL  FILL_4020
timestamp 1018054153
transform 1 0 6432 0 1 5280
box -16 -6 32 210
use FILL  FILL_4022
timestamp 1018054153
transform 1 0 6448 0 1 5280
box -16 -6 32 210
use FILL  FILL_4023
timestamp 1018054153
transform 1 0 6464 0 1 5280
box -16 -6 32 210
use FILL  FILL_4024
timestamp 1018054153
transform 1 0 6480 0 1 5280
box -16 -6 32 210
use FILL  FILL_4025
timestamp 1018054153
transform 1 0 6496 0 1 5280
box -16 -6 32 210
use FILL  FILL_4026
timestamp 1018054153
transform 1 0 6512 0 1 5280
box -16 -6 32 210
use FILL  FILL_4027
timestamp 1018054153
transform 1 0 6528 0 1 5280
box -16 -6 32 210
use FILL  FILL_4030
timestamp 1018054153
transform 1 0 6544 0 1 5280
box -16 -6 32 210
use FILL  FILL_4032
timestamp 1018054153
transform 1 0 6560 0 1 5280
box -16 -6 32 210
use FILL  FILL_4034
timestamp 1018054153
transform 1 0 6576 0 1 5280
box -16 -6 32 210
use FILL  FILL_4036
timestamp 1018054153
transform 1 0 6592 0 1 5280
box -16 -6 32 210
use FILL  FILL_4038
timestamp 1018054153
transform 1 0 6608 0 1 5280
box -16 -6 32 210
use FILL  FILL_4040
timestamp 1018054153
transform 1 0 6624 0 1 5280
box -16 -6 32 210
use FILL  FILL_4042
timestamp 1018054153
transform 1 0 6640 0 1 5280
box -16 -6 32 210
use FILL  FILL_4044
timestamp 1018054153
transform 1 0 6656 0 1 5280
box -16 -6 32 210
use FILL  FILL_4046
timestamp 1018054153
transform 1 0 6672 0 1 5280
box -16 -6 32 210
use FILL  FILL_4048
timestamp 1018054153
transform 1 0 6688 0 1 5280
box -16 -6 32 210
use FILL  FILL_4050
timestamp 1018054153
transform 1 0 6704 0 1 5280
box -16 -6 32 210
use FILL  FILL_4052
timestamp 1018054153
transform 1 0 6720 0 1 5280
box -16 -6 32 210
use FILL  FILL_4054
timestamp 1018054153
transform 1 0 6736 0 1 5280
box -16 -6 32 210
use FILL  FILL_4056
timestamp 1018054153
transform 1 0 6752 0 1 5280
box -16 -6 32 210
use AND2X2  AND2X2_1
timestamp 1090541974
transform 1 0 6768 0 1 5280
box -16 -6 80 210
use FILL  FILL_4058
timestamp 1018054153
transform 1 0 6832 0 1 5280
box -16 -6 32 210
use FILL  FILL_4064
timestamp 1018054153
transform 1 0 6848 0 1 5280
box -16 -6 32 210
use FILL  FILL_4066
timestamp 1018054153
transform 1 0 6864 0 1 5280
box -16 -6 32 210
use FILL  FILL_4068
timestamp 1018054153
transform 1 0 6880 0 1 5280
box -16 -6 32 210
use FILL  FILL_4070
timestamp 1018054153
transform 1 0 6896 0 1 5280
box -16 -6 32 210
use FILL  FILL_4072
timestamp 1018054153
transform 1 0 6912 0 1 5280
box -16 -6 32 210
use FILL  FILL_4074
timestamp 1018054153
transform 1 0 6928 0 1 5280
box -16 -6 32 210
use FILL  FILL_4076
timestamp 1018054153
transform 1 0 6944 0 1 5280
box -16 -6 32 210
use FILL  FILL_4078
timestamp 1018054153
transform 1 0 6960 0 1 5280
box -16 -6 32 210
use FILL  FILL_4080
timestamp 1018054153
transform 1 0 6976 0 1 5280
box -16 -6 32 210
use FILL  FILL_4082
timestamp 1018054153
transform 1 0 6992 0 1 5280
box -16 -6 32 210
use FILL  FILL_4084
timestamp 1018054153
transform 1 0 7008 0 1 5280
box -16 -6 32 210
use FILL  FILL_4086
timestamp 1018054153
transform 1 0 7024 0 1 5280
box -16 -6 32 210
use FILL  FILL_4088
timestamp 1018054153
transform 1 0 7040 0 1 5280
box -16 -6 32 210
use FILL  FILL_4090
timestamp 1018054153
transform 1 0 7056 0 1 5280
box -16 -6 32 210
use FILL  FILL_4092
timestamp 1018054153
transform 1 0 7072 0 1 5280
box -16 -6 32 210
use FILL  FILL_4094
timestamp 1018054153
transform 1 0 7088 0 1 5280
box -16 -6 32 210
use FILL  FILL_4096
timestamp 1018054153
transform 1 0 7104 0 1 5280
box -16 -6 32 210
use FILL  FILL_4098
timestamp 1018054153
transform 1 0 7120 0 1 5280
box -16 -6 32 210
use FILL  FILL_4100
timestamp 1018054153
transform 1 0 7136 0 1 5280
box -16 -6 32 210
use FILL  FILL_4102
timestamp 1018054153
transform 1 0 7152 0 1 5280
box -16 -6 32 210
use FILL  FILL_4104
timestamp 1018054153
transform 1 0 7168 0 1 5280
box -16 -6 32 210
use FILL  FILL_4106
timestamp 1018054153
transform 1 0 7184 0 1 5280
box -16 -6 32 210
use FILL  FILL_4108
timestamp 1018054153
transform 1 0 7200 0 1 5280
box -16 -6 32 210
use FILL  FILL_4110
timestamp 1018054153
transform 1 0 7216 0 1 5280
box -16 -6 32 210
use FILL  FILL_4112
timestamp 1018054153
transform 1 0 7232 0 1 5280
box -16 -6 32 210
use FILL  FILL_4114
timestamp 1018054153
transform 1 0 7248 0 1 5280
box -16 -6 32 210
use FILL  FILL_4116
timestamp 1018054153
transform 1 0 7264 0 1 5280
box -16 -6 32 210
use FILL  FILL_4118
timestamp 1018054153
transform 1 0 7280 0 1 5280
box -16 -6 32 210
use FILL  FILL_4120
timestamp 1018054153
transform 1 0 7296 0 1 5280
box -16 -6 32 210
use FILL  FILL_4122
timestamp 1018054153
transform 1 0 7312 0 1 5280
box -16 -6 32 210
use FILL  FILL_4124
timestamp 1018054153
transform 1 0 7328 0 1 5280
box -16 -6 32 210
use FILL  FILL_4126
timestamp 1018054153
transform 1 0 7344 0 1 5280
box -16 -6 32 210
use FILL  FILL_4128
timestamp 1018054153
transform 1 0 7360 0 1 5280
box -16 -6 32 210
use FILL  FILL_4130
timestamp 1018054153
transform 1 0 7376 0 1 5280
box -16 -6 32 210
use FILL  FILL_4132
timestamp 1018054153
transform 1 0 7392 0 1 5280
box -16 -6 32 210
use FILL  FILL_4134
timestamp 1018054153
transform 1 0 7408 0 1 5280
box -16 -6 32 210
use FILL  FILL_4136
timestamp 1018054153
transform 1 0 7424 0 1 5280
box -16 -6 32 210
use FILL  FILL_4138
timestamp 1018054153
transform 1 0 7440 0 1 5280
box -16 -6 32 210
use FILL  FILL_4140
timestamp 1018054153
transform 1 0 7456 0 1 5280
box -16 -6 32 210
use FILL  FILL_4142
timestamp 1018054153
transform 1 0 7472 0 1 5280
box -16 -6 32 210
use FILL  FILL_4144
timestamp 1018054153
transform 1 0 7488 0 1 5280
box -16 -6 32 210
use FILL  FILL_4146
timestamp 1018054153
transform 1 0 7504 0 1 5280
box -16 -6 32 210
use FILL  FILL_4148
timestamp 1018054153
transform 1 0 7520 0 1 5280
box -16 -6 32 210
use FILL  FILL_4150
timestamp 1018054153
transform 1 0 7536 0 1 5280
box -16 -6 32 210
use FILL  FILL_4152
timestamp 1018054153
transform 1 0 7552 0 1 5280
box -16 -6 32 210
use FILL  FILL_4154
timestamp 1018054153
transform 1 0 7568 0 1 5280
box -16 -6 32 210
use FILL  FILL_4156
timestamp 1018054153
transform 1 0 7584 0 1 5280
box -16 -6 32 210
use FILL  FILL_4158
timestamp 1018054153
transform 1 0 7600 0 1 5280
box -16 -6 32 210
use FILL  FILL_4160
timestamp 1018054153
transform 1 0 7616 0 1 5280
box -16 -6 32 210
use FILL  FILL_4162
timestamp 1018054153
transform 1 0 7632 0 1 5280
box -16 -6 32 210
use FILL  FILL_4164
timestamp 1018054153
transform 1 0 7648 0 1 5280
box -16 -6 32 210
use FILL  FILL_4166
timestamp 1018054153
transform 1 0 7664 0 1 5280
box -16 -6 32 210
use FILL  FILL_4168
timestamp 1018054153
transform 1 0 7680 0 1 5280
box -16 -6 32 210
use FILL  FILL_4170
timestamp 1018054153
transform 1 0 7696 0 1 5280
box -16 -6 32 210
use FILL  FILL_4172
timestamp 1018054153
transform 1 0 7712 0 1 5280
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_21
timestamp 1542725905
transform 1 0 7908 0 1 5280
box -48 -6 48 6
use M3_M2  M3_M2_65
timestamp 1542725905
transform 1 0 3528 0 1 5210
box -6 -6 6 6
use M2_M1  M2_M1_181
timestamp 1542725905
transform 1 0 4392 0 1 5230
box -4 -4 4 4
use M2_M1  M2_M1_184
timestamp 1542725905
transform 1 0 4488 0 1 5210
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_22
timestamp 1542725905
transform 1 0 2212 0 1 5080
box -48 -6 48 6
use PADINC  PADINC_6
timestamp 1084294328
transform 0 -1 2000 1 0 5000
box -12 -6 606 2000
use M3_M2  M3_M2_73
timestamp 1542725905
transform 1 0 1998 0 1 4930
box -6 -6 6 6
use FILL  FILL_3549
timestamp 1018054153
transform 1 0 2272 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3551
timestamp 1018054153
transform 1 0 2288 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3553
timestamp 1018054153
transform 1 0 2304 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3555
timestamp 1018054153
transform 1 0 2320 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3557
timestamp 1018054153
transform 1 0 2336 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3559
timestamp 1018054153
transform 1 0 2352 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3561
timestamp 1018054153
transform 1 0 2368 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3563
timestamp 1018054153
transform 1 0 2384 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3565
timestamp 1018054153
transform 1 0 2400 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3567
timestamp 1018054153
transform 1 0 2416 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3569
timestamp 1018054153
transform 1 0 2432 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3571
timestamp 1018054153
transform 1 0 2448 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3573
timestamp 1018054153
transform 1 0 2464 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3575
timestamp 1018054153
transform 1 0 2480 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3577
timestamp 1018054153
transform 1 0 2496 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3579
timestamp 1018054153
transform 1 0 2512 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3581
timestamp 1018054153
transform 1 0 2528 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3583
timestamp 1018054153
transform 1 0 2544 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3585
timestamp 1018054153
transform 1 0 2560 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3587
timestamp 1018054153
transform 1 0 2576 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3589
timestamp 1018054153
transform 1 0 2592 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3591
timestamp 1018054153
transform 1 0 2608 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3593
timestamp 1018054153
transform 1 0 2624 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3595
timestamp 1018054153
transform 1 0 2640 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3597
timestamp 1018054153
transform 1 0 2656 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3599
timestamp 1018054153
transform 1 0 2672 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3601
timestamp 1018054153
transform 1 0 2688 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3603
timestamp 1018054153
transform 1 0 2704 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3605
timestamp 1018054153
transform 1 0 2720 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3607
timestamp 1018054153
transform 1 0 2736 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3609
timestamp 1018054153
transform 1 0 2752 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3611
timestamp 1018054153
transform 1 0 2768 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3613
timestamp 1018054153
transform 1 0 2784 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3615
timestamp 1018054153
transform 1 0 2800 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3617
timestamp 1018054153
transform 1 0 2816 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3619
timestamp 1018054153
transform 1 0 2832 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3621
timestamp 1018054153
transform 1 0 2848 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3623
timestamp 1018054153
transform 1 0 2864 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3625
timestamp 1018054153
transform 1 0 2880 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3627
timestamp 1018054153
transform 1 0 2896 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3629
timestamp 1018054153
transform 1 0 2912 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3631
timestamp 1018054153
transform 1 0 2928 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3633
timestamp 1018054153
transform 1 0 2944 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3635
timestamp 1018054153
transform 1 0 2960 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3637
timestamp 1018054153
transform 1 0 2976 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3639
timestamp 1018054153
transform 1 0 2992 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3641
timestamp 1018054153
transform 1 0 3008 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3643
timestamp 1018054153
transform 1 0 3024 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3645
timestamp 1018054153
transform 1 0 3040 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3647
timestamp 1018054153
transform 1 0 3056 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3649
timestamp 1018054153
transform 1 0 3072 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3651
timestamp 1018054153
transform 1 0 3088 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3653
timestamp 1018054153
transform 1 0 3104 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3655
timestamp 1018054153
transform 1 0 3120 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3657
timestamp 1018054153
transform 1 0 3136 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3659
timestamp 1018054153
transform 1 0 3152 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3661
timestamp 1018054153
transform 1 0 3168 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3663
timestamp 1018054153
transform 1 0 3184 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3665
timestamp 1018054153
transform 1 0 3200 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3667
timestamp 1018054153
transform 1 0 3216 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3669
timestamp 1018054153
transform 1 0 3232 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3671
timestamp 1018054153
transform 1 0 3248 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3673
timestamp 1018054153
transform 1 0 3264 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3675
timestamp 1018054153
transform 1 0 3280 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3677
timestamp 1018054153
transform 1 0 3296 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3679
timestamp 1018054153
transform 1 0 3312 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3681
timestamp 1018054153
transform 1 0 3328 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3683
timestamp 1018054153
transform 1 0 3344 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3685
timestamp 1018054153
transform 1 0 3360 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3687
timestamp 1018054153
transform 1 0 3376 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3689
timestamp 1018054153
transform 1 0 3392 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3691
timestamp 1018054153
transform 1 0 3408 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3693
timestamp 1018054153
transform 1 0 3424 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3695
timestamp 1018054153
transform 1 0 3440 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3697
timestamp 1018054153
transform 1 0 3456 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3699
timestamp 1018054153
transform 1 0 3472 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3701
timestamp 1018054153
transform 1 0 3488 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3703
timestamp 1018054153
transform 1 0 3504 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3705
timestamp 1018054153
transform 1 0 3520 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3707
timestamp 1018054153
transform 1 0 3536 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3709
timestamp 1018054153
transform 1 0 3552 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3711
timestamp 1018054153
transform 1 0 3568 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3713
timestamp 1018054153
transform 1 0 3584 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3715
timestamp 1018054153
transform 1 0 3600 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3717
timestamp 1018054153
transform 1 0 3616 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3719
timestamp 1018054153
transform 1 0 3632 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3721
timestamp 1018054153
transform 1 0 3648 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3723
timestamp 1018054153
transform 1 0 3664 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3725
timestamp 1018054153
transform 1 0 3680 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3727
timestamp 1018054153
transform 1 0 3696 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3729
timestamp 1018054153
transform 1 0 3712 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3731
timestamp 1018054153
transform 1 0 3728 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3733
timestamp 1018054153
transform 1 0 3744 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3735
timestamp 1018054153
transform 1 0 3760 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3737
timestamp 1018054153
transform 1 0 3776 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3739
timestamp 1018054153
transform 1 0 3792 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3741
timestamp 1018054153
transform 1 0 3808 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3743
timestamp 1018054153
transform 1 0 3824 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3745
timestamp 1018054153
transform 1 0 3840 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3747
timestamp 1018054153
transform 1 0 3856 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3749
timestamp 1018054153
transform 1 0 3872 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3751
timestamp 1018054153
transform 1 0 3888 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3753
timestamp 1018054153
transform 1 0 3904 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3755
timestamp 1018054153
transform 1 0 3920 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3757
timestamp 1018054153
transform 1 0 3936 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3759
timestamp 1018054153
transform 1 0 3952 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3761
timestamp 1018054153
transform 1 0 3968 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3763
timestamp 1018054153
transform 1 0 3984 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3765
timestamp 1018054153
transform 1 0 4000 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3767
timestamp 1018054153
transform 1 0 4016 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3769
timestamp 1018054153
transform 1 0 4032 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3771
timestamp 1018054153
transform 1 0 4048 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3773
timestamp 1018054153
transform 1 0 4064 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3775
timestamp 1018054153
transform 1 0 4080 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3777
timestamp 1018054153
transform 1 0 4096 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3779
timestamp 1018054153
transform 1 0 4112 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3781
timestamp 1018054153
transform 1 0 4128 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3783
timestamp 1018054153
transform 1 0 4144 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3785
timestamp 1018054153
transform 1 0 4160 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3787
timestamp 1018054153
transform 1 0 4176 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3789
timestamp 1018054153
transform 1 0 4192 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3791
timestamp 1018054153
transform 1 0 4208 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3792
timestamp 1018054153
transform 1 0 4224 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3793
timestamp 1018054153
transform 1 0 4240 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3795
timestamp 1018054153
transform 1 0 4256 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3797
timestamp 1018054153
transform 1 0 4272 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3799
timestamp 1018054153
transform 1 0 4288 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3801
timestamp 1018054153
transform 1 0 4304 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3803
timestamp 1018054153
transform 1 0 4320 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3805
timestamp 1018054153
transform 1 0 4336 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3807
timestamp 1018054153
transform 1 0 4352 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3809
timestamp 1018054153
transform 1 0 4368 0 -1 5280
box -16 -6 32 210
use INVX1  INVX1_10
timestamp 1053022145
transform 1 0 4384 0 -1 5280
box -18 -6 52 210
use FILL  FILL_3813
timestamp 1018054153
transform 1 0 4416 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3815
timestamp 1018054153
transform 1 0 4432 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3817
timestamp 1018054153
transform 1 0 4448 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3819
timestamp 1018054153
transform 1 0 4464 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3821
timestamp 1018054153
transform 1 0 4480 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3823
timestamp 1018054153
transform 1 0 4496 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3824
timestamp 1018054153
transform 1 0 4512 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3825
timestamp 1018054153
transform 1 0 4528 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3826
timestamp 1018054153
transform 1 0 4544 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3828
timestamp 1018054153
transform 1 0 4560 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3830
timestamp 1018054153
transform 1 0 4576 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3832
timestamp 1018054153
transform 1 0 4592 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3834
timestamp 1018054153
transform 1 0 4608 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3836
timestamp 1018054153
transform 1 0 4624 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_194
timestamp 1542725905
transform 1 0 4664 0 1 5190
box -4 -4 4 4
use FILL  FILL_3838
timestamp 1018054153
transform 1 0 4640 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3840
timestamp 1018054153
transform 1 0 4656 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_185
timestamp 1542725905
transform 1 0 4696 0 1 5210
box -4 -4 4 4
use FILL  FILL_3842
timestamp 1018054153
transform 1 0 4672 0 -1 5280
box -16 -6 32 210
use OAI21X1  OAI21X1_11
timestamp 1053722159
transform 1 0 4688 0 -1 5280
box -16 -6 68 210
use M2_M1  M2_M1_186
timestamp 1542725905
transform 1 0 4760 0 1 5210
box -4 -4 4 4
use FILL  FILL_3848
timestamp 1018054153
transform 1 0 4752 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3849
timestamp 1018054153
transform 1 0 4768 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3850
timestamp 1018054153
transform 1 0 4784 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3851
timestamp 1018054153
transform 1 0 4800 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3853
timestamp 1018054153
transform 1 0 4816 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3855
timestamp 1018054153
transform 1 0 4832 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3857
timestamp 1018054153
transform 1 0 4848 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3859
timestamp 1018054153
transform 1 0 4864 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3861
timestamp 1018054153
transform 1 0 4880 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3863
timestamp 1018054153
transform 1 0 4896 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3865
timestamp 1018054153
transform 1 0 4912 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3867
timestamp 1018054153
transform 1 0 4928 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_187
timestamp 1542725905
transform 1 0 4968 0 1 5210
box -4 -4 4 4
use FILL  FILL_3869
timestamp 1018054153
transform 1 0 4944 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3871
timestamp 1018054153
transform 1 0 4960 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3877
timestamp 1018054153
transform 1 0 4976 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_188
timestamp 1542725905
transform 1 0 5096 0 1 5210
box -4 -4 4 4
use M2_M1  M2_M1_195
timestamp 1542725905
transform 1 0 5048 0 1 5190
box -4 -4 4 4
use XOR2X1  XOR2X1_3
timestamp 1053359338
transform -1 0 5104 0 -1 5280
box -16 -6 128 210
use FILL  FILL_3878
timestamp 1018054153
transform 1 0 5104 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3880
timestamp 1018054153
transform 1 0 5120 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3882
timestamp 1018054153
transform 1 0 5136 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3884
timestamp 1018054153
transform 1 0 5152 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3886
timestamp 1018054153
transform 1 0 5168 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3888
timestamp 1018054153
transform 1 0 5184 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3890
timestamp 1018054153
transform 1 0 5200 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3892
timestamp 1018054153
transform 1 0 5216 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3894
timestamp 1018054153
transform 1 0 5232 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3896
timestamp 1018054153
transform 1 0 5248 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3898
timestamp 1018054153
transform 1 0 5264 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3900
timestamp 1018054153
transform 1 0 5280 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3901
timestamp 1018054153
transform 1 0 5296 0 -1 5280
box -16 -6 32 210
use M3_M2  M3_M2_64
timestamp 1542725905
transform 1 0 5336 0 1 5250
box -6 -6 6 6
use M2_M1  M2_M1_182
timestamp 1542725905
transform 1 0 5336 0 1 5230
box -4 -4 4 4
use FILL  FILL_3902
timestamp 1018054153
transform 1 0 5312 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_189
timestamp 1542725905
transform 1 0 5368 0 1 5210
box -4 -4 4 4
use INVX1  INVX1_12
timestamp 1053022145
transform 1 0 5328 0 -1 5280
box -18 -6 52 210
use FILL  FILL_3906
timestamp 1018054153
transform 1 0 5360 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3908
timestamp 1018054153
transform 1 0 5376 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3910
timestamp 1018054153
transform 1 0 5392 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3912
timestamp 1018054153
transform 1 0 5408 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3914
timestamp 1018054153
transform 1 0 5424 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3916
timestamp 1018054153
transform 1 0 5440 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3918
timestamp 1018054153
transform 1 0 5456 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_190
timestamp 1542725905
transform 1 0 5496 0 1 5210
box -4 -4 4 4
use FILL  FILL_3920
timestamp 1018054153
transform 1 0 5472 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3922
timestamp 1018054153
transform 1 0 5488 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3924
timestamp 1018054153
transform 1 0 5504 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3925
timestamp 1018054153
transform 1 0 5520 0 -1 5280
box -16 -6 32 210
use M3_M2  M3_M2_66
timestamp 1542725905
transform 1 0 5560 0 1 5150
box -6 -6 6 6
use FILL  FILL_3926
timestamp 1018054153
transform 1 0 5536 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3927
timestamp 1018054153
transform 1 0 5552 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3929
timestamp 1018054153
transform 1 0 5568 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3931
timestamp 1018054153
transform 1 0 5584 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3933
timestamp 1018054153
transform 1 0 5600 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3935
timestamp 1018054153
transform 1 0 5616 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3937
timestamp 1018054153
transform 1 0 5632 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3939
timestamp 1018054153
transform 1 0 5648 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3941
timestamp 1018054153
transform 1 0 5664 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3943
timestamp 1018054153
transform 1 0 5680 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3945
timestamp 1018054153
transform 1 0 5696 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3947
timestamp 1018054153
transform 1 0 5712 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3949
timestamp 1018054153
transform 1 0 5728 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3951
timestamp 1018054153
transform 1 0 5744 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3952
timestamp 1018054153
transform 1 0 5760 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3953
timestamp 1018054153
transform 1 0 5776 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3955
timestamp 1018054153
transform 1 0 5792 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3957
timestamp 1018054153
transform 1 0 5808 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3959
timestamp 1018054153
transform 1 0 5824 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_191
timestamp 1542725905
transform 1 0 5864 0 1 5210
box -4 -4 4 4
use FILL  FILL_3961
timestamp 1018054153
transform 1 0 5840 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3963
timestamp 1018054153
transform 1 0 5856 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3965
timestamp 1018054153
transform 1 0 5872 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3967
timestamp 1018054153
transform 1 0 5888 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3969
timestamp 1018054153
transform 1 0 5904 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_192
timestamp 1542725905
transform 1 0 6024 0 1 5210
box -4 -4 4 4
use M2_M1  M2_M1_196
timestamp 1542725905
transform 1 0 5976 0 1 5190
box -4 -4 4 4
use XOR2X1  XOR2X1_4
timestamp 1053359338
transform 1 0 5920 0 -1 5280
box -16 -6 128 210
use FILL  FILL_3978
timestamp 1018054153
transform 1 0 6032 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3980
timestamp 1018054153
transform 1 0 6048 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3982
timestamp 1018054153
transform 1 0 6064 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3984
timestamp 1018054153
transform 1 0 6080 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3986
timestamp 1018054153
transform 1 0 6096 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3988
timestamp 1018054153
transform 1 0 6112 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3990
timestamp 1018054153
transform 1 0 6128 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3992
timestamp 1018054153
transform 1 0 6144 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3994
timestamp 1018054153
transform 1 0 6160 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3996
timestamp 1018054153
transform 1 0 6176 0 -1 5280
box -16 -6 32 210
use FILL  FILL_3998
timestamp 1018054153
transform 1 0 6192 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4000
timestamp 1018054153
transform 1 0 6208 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4002
timestamp 1018054153
transform 1 0 6224 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4004
timestamp 1018054153
transform 1 0 6240 0 -1 5280
box -16 -6 32 210
use M3_M2  M3_M2_67
timestamp 1542725905
transform 1 0 6280 0 1 5150
box -6 -6 6 6
use FILL  FILL_4006
timestamp 1018054153
transform 1 0 6256 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4008
timestamp 1018054153
transform 1 0 6272 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4009
timestamp 1018054153
transform 1 0 6288 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4010
timestamp 1018054153
transform 1 0 6304 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4011
timestamp 1018054153
transform 1 0 6320 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4012
timestamp 1018054153
transform 1 0 6336 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4013
timestamp 1018054153
transform 1 0 6352 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4014
timestamp 1018054153
transform 1 0 6368 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4015
timestamp 1018054153
transform 1 0 6384 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4017
timestamp 1018054153
transform 1 0 6400 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_197
timestamp 1542725905
transform 1 0 6440 0 1 5190
box -4 -4 4 4
use FILL  FILL_4019
timestamp 1018054153
transform 1 0 6416 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4021
timestamp 1018054153
transform 1 0 6432 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4028
timestamp 1018054153
transform 1 0 6448 0 -1 5280
box -16 -6 32 210
use OR2X1  OR2X1_0
timestamp 1090542464
transform -1 0 6528 0 -1 5280
box -16 -6 80 210
use FILL  FILL_4029
timestamp 1018054153
transform 1 0 6528 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_183
timestamp 1542725905
transform 1 0 6568 0 1 5230
box -4 -4 4 4
use FILL  FILL_4031
timestamp 1018054153
transform 1 0 6544 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_193
timestamp 1542725905
transform 1 0 6824 0 1 5210
box -4 -4 4 4
use FILL  FILL_4033
timestamp 1018054153
transform 1 0 6560 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4035
timestamp 1018054153
transform 1 0 6576 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4037
timestamp 1018054153
transform 1 0 6592 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4039
timestamp 1018054153
transform 1 0 6608 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4041
timestamp 1018054153
transform 1 0 6624 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4043
timestamp 1018054153
transform 1 0 6640 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4045
timestamp 1018054153
transform 1 0 6656 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4047
timestamp 1018054153
transform 1 0 6672 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4049
timestamp 1018054153
transform 1 0 6688 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4051
timestamp 1018054153
transform 1 0 6704 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4053
timestamp 1018054153
transform 1 0 6720 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4055
timestamp 1018054153
transform 1 0 6736 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4057
timestamp 1018054153
transform 1 0 6752 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4059
timestamp 1018054153
transform 1 0 6768 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4060
timestamp 1018054153
transform 1 0 6784 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4061
timestamp 1018054153
transform 1 0 6800 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4062
timestamp 1018054153
transform 1 0 6816 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4063
timestamp 1018054153
transform 1 0 6832 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4065
timestamp 1018054153
transform 1 0 6848 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4067
timestamp 1018054153
transform 1 0 6864 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4069
timestamp 1018054153
transform 1 0 6880 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4071
timestamp 1018054153
transform 1 0 6896 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4073
timestamp 1018054153
transform 1 0 6912 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4075
timestamp 1018054153
transform 1 0 6928 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4077
timestamp 1018054153
transform 1 0 6944 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4079
timestamp 1018054153
transform 1 0 6960 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4081
timestamp 1018054153
transform 1 0 6976 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4083
timestamp 1018054153
transform 1 0 6992 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4085
timestamp 1018054153
transform 1 0 7008 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4087
timestamp 1018054153
transform 1 0 7024 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4089
timestamp 1018054153
transform 1 0 7040 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4091
timestamp 1018054153
transform 1 0 7056 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4093
timestamp 1018054153
transform 1 0 7072 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4095
timestamp 1018054153
transform 1 0 7088 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4097
timestamp 1018054153
transform 1 0 7104 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4099
timestamp 1018054153
transform 1 0 7120 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4101
timestamp 1018054153
transform 1 0 7136 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4103
timestamp 1018054153
transform 1 0 7152 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4105
timestamp 1018054153
transform 1 0 7168 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4107
timestamp 1018054153
transform 1 0 7184 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4109
timestamp 1018054153
transform 1 0 7200 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4111
timestamp 1018054153
transform 1 0 7216 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4113
timestamp 1018054153
transform 1 0 7232 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4115
timestamp 1018054153
transform 1 0 7248 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4117
timestamp 1018054153
transform 1 0 7264 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4119
timestamp 1018054153
transform 1 0 7280 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4121
timestamp 1018054153
transform 1 0 7296 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4123
timestamp 1018054153
transform 1 0 7312 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4125
timestamp 1018054153
transform 1 0 7328 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4127
timestamp 1018054153
transform 1 0 7344 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4129
timestamp 1018054153
transform 1 0 7360 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4131
timestamp 1018054153
transform 1 0 7376 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4133
timestamp 1018054153
transform 1 0 7392 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4135
timestamp 1018054153
transform 1 0 7408 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4137
timestamp 1018054153
transform 1 0 7424 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4139
timestamp 1018054153
transform 1 0 7440 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4141
timestamp 1018054153
transform 1 0 7456 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4143
timestamp 1018054153
transform 1 0 7472 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4145
timestamp 1018054153
transform 1 0 7488 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4147
timestamp 1018054153
transform 1 0 7504 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4149
timestamp 1018054153
transform 1 0 7520 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4151
timestamp 1018054153
transform 1 0 7536 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4153
timestamp 1018054153
transform 1 0 7552 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4155
timestamp 1018054153
transform 1 0 7568 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4157
timestamp 1018054153
transform 1 0 7584 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4159
timestamp 1018054153
transform 1 0 7600 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4161
timestamp 1018054153
transform 1 0 7616 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4163
timestamp 1018054153
transform 1 0 7632 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4165
timestamp 1018054153
transform 1 0 7648 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4167
timestamp 1018054153
transform 1 0 7664 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4169
timestamp 1018054153
transform 1 0 7680 0 -1 5280
box -16 -6 32 210
use FILL  FILL_4171
timestamp 1018054153
transform 1 0 7696 0 -1 5280
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_23
timestamp 1542725905
transform 1 0 7788 0 1 5080
box -48 -6 48 6
use FILL  FILL_4173
timestamp 1018054153
transform 1 0 7712 0 -1 5280
box -16 -6 32 210
use M2_M1  M2_M1_212
timestamp 1542725905
transform 1 0 3800 0 1 4950
box -4 -4 4 4
use M2_M1  M2_M1_201
timestamp 1542725905
transform 1 0 3848 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_202
timestamp 1542725905
transform 1 0 4120 0 1 4970
box -4 -4 4 4
use M3_M2  M3_M2_75
timestamp 1542725905
transform 1 0 4392 0 1 4910
box -6 -6 6 6
use M3_M2  M3_M2_70
timestamp 1542725905
transform 1 0 4456 0 1 4990
box -6 -6 6 6
use M2_M1  M2_M1_213
timestamp 1542725905
transform 1 0 4456 0 1 4950
box -4 -4 4 4
use M2_M1  M2_M1_203
timestamp 1542725905
transform 1 0 4488 0 1 4970
box -4 -4 4 4
use mult_pad_VIA2  mult_pad_VIA2_0
timestamp 1542725905
transform 1 0 4625 0 1 5031
box -6 -6 6 6
use mult_pad_VIA3  mult_pad_VIA3_0
timestamp 1542725905
transform 1 0 4709 0 1 5031
box -10 -6 10 6
use M2_M1  M2_M1_198
timestamp 1542725905
transform 1 0 4824 0 1 5030
box -4 -4 4 4
use mult_pad_VIA7  mult_pad_VIA7_0
timestamp 1542725905
transform 1 0 5147 0 1 5031
box -20 -6 20 6
use mult_pad_VIA7  mult_pad_VIA7_1
timestamp 1542725905
transform 1 0 5595 0 1 5031
box -20 -6 20 6
use mult_pad_VIA7  mult_pad_VIA7_2
timestamp 1542725905
transform 1 0 6043 0 1 5031
box -20 -6 20 6
use M3_M2  M3_M2_68
timestamp 1542725905
transform 1 0 6408 0 1 5030
box -6 -6 6 6
use mult_pad_VIA3  mult_pad_VIA3_1
timestamp 1542725905
transform 1 0 6481 0 1 5031
box -10 -6 10 6
use mult_pad_VIA2  mult_pad_VIA2_1
timestamp 1542725905
transform 1 0 6565 0 1 5031
box -6 -6 6 6
use mult_pad_VIA2  mult_pad_VIA2_2
timestamp 1542725905
transform 1 0 4649 0 1 5007
box -6 -6 6 6
use mult_pad_VIA12  mult_pad_VIA12_0
timestamp 1542725905
transform 1 0 4923 0 1 5007
box -16 -6 16 6
use mult_pad_VIA12  mult_pad_VIA12_1
timestamp 1542725905
transform 1 0 5371 0 1 5007
box -16 -6 16 6
use M3_M2  M3_M2_69
timestamp 1542725905
transform 1 0 5512 0 1 5010
box -6 -6 6 6
use mult_pad_VIA12  mult_pad_VIA12_2
timestamp 1542725905
transform 1 0 5819 0 1 5007
box -16 -6 16 6
use mult_pad_VIA12  mult_pad_VIA12_3
timestamp 1542725905
transform 1 0 6267 0 1 5007
box -16 -6 16 6
use mult_pad_VIA2  mult_pad_VIA2_3
timestamp 1542725905
transform 1 0 6541 0 1 5007
box -6 -6 6 6
use M3_M2  M3_M2_71
timestamp 1542725905
transform 1 0 5016 0 1 4990
box -6 -6 6 6
use M2_M1  M2_M1_199
timestamp 1542725905
transform 1 0 5736 0 1 4990
box -4 -4 4 4
use M2_M1  M2_M1_204
timestamp 1542725905
transform 1 0 4888 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_205
timestamp 1542725905
transform 1 0 5016 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_206
timestamp 1542725905
transform 1 0 5208 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_207
timestamp 1542725905
transform 1 0 5320 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_208
timestamp 1542725905
transform 1 0 5656 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_209
timestamp 1542725905
transform 1 0 5752 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_210
timestamp 1542725905
transform 1 0 5896 0 1 4970
box -4 -4 4 4
use mult_pad_VIA4  mult_pad_VIA4_0
timestamp 1542725905
transform 1 0 4709 0 1 4947
box -10 -10 10 10
use M2_M1  M2_M1_214
timestamp 1542725905
transform 1 0 4783 0 1 4950
box -4 -4 4 4
use M2_M1  M2_M1_215
timestamp 1542725905
transform 1 0 4824 0 1 4950
box -4 -4 4 4
use mult_pad_VIA9  mult_pad_VIA9_0
timestamp 1542725905
transform 1 0 4923 0 1 4957
box -16 -4 16 4
use mult_pad_VIA8  mult_pad_VIA8_0
timestamp 1542725905
transform 1 0 4923 0 1 4953
box -4 -4 4 4
use M2_M1  M2_M1_216
timestamp 1542725905
transform 1 0 5064 0 1 4950
box -4 -4 4 4
use mult_pad_VIA5  mult_pad_VIA5_0
timestamp 1542725905
transform 1 0 5147 0 1 4955
box -20 -4 20 4
use mult_pad_VIA11  mult_pad_VIA11_0
timestamp 1542725905
transform 1 0 5371 0 1 4955
box -16 -4 16 4
use M2_M1  M2_M1_217
timestamp 1542725905
transform 1 0 5512 0 1 4950
box -4 -4 4 4
use mult_pad_VIA5  mult_pad_VIA5_1
timestamp 1542725905
transform 1 0 5595 0 1 4955
box -20 -4 20 4
use M3_M2  M3_M2_72
timestamp 1542725905
transform 1 0 5752 0 1 4950
box -6 -6 6 6
use mult_pad_VIA11  mult_pad_VIA11_1
timestamp 1542725905
transform 1 0 5819 0 1 4955
box -16 -4 16 4
use M2_M1  M2_M1_218
timestamp 1542725905
transform 1 0 5960 0 1 4950
box -4 -4 4 4
use mult_pad_VIA5  mult_pad_VIA5_2
timestamp 1542725905
transform 1 0 6043 0 1 4955
box -20 -4 20 4
use M2_M1  M2_M1_219
timestamp 1542725905
transform 1 0 6127 0 1 4950
box -4 -4 4 4
use mult_pad_VIA9  mult_pad_VIA9_1
timestamp 1542725905
transform 1 0 6267 0 1 4955
box -16 -4 16 4
use mult_pad_VIA8  mult_pad_VIA8_1
timestamp 1542725905
transform 1 0 6267 0 1 4953
box -4 -4 4 4
use M2_M1  M2_M1_220
timestamp 1542725905
transform 1 0 6408 0 1 4950
box -4 -4 4 4
use mult_pad_VIA4  mult_pad_VIA4_1
timestamp 1542725905
transform 1 0 6481 0 1 4947
box -10 -10 10 10
use M3_M2  M3_M2_74
timestamp 1542725905
transform 1 0 5896 0 1 4930
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_24
timestamp 1542725905
transform 1 0 2092 0 1 4880
box -48 -6 48 6
use FILL  FILL_4174
timestamp 1018054153
transform 1 0 2272 0 1 4880
box -16 -6 32 210
use FILL  FILL_4176
timestamp 1018054153
transform 1 0 2288 0 1 4880
box -16 -6 32 210
use FILL  FILL_4178
timestamp 1018054153
transform 1 0 2304 0 1 4880
box -16 -6 32 210
use FILL  FILL_4180
timestamp 1018054153
transform 1 0 2320 0 1 4880
box -16 -6 32 210
use FILL  FILL_4182
timestamp 1018054153
transform 1 0 2336 0 1 4880
box -16 -6 32 210
use FILL  FILL_4184
timestamp 1018054153
transform 1 0 2352 0 1 4880
box -16 -6 32 210
use FILL  FILL_4186
timestamp 1018054153
transform 1 0 2368 0 1 4880
box -16 -6 32 210
use FILL  FILL_4188
timestamp 1018054153
transform 1 0 2384 0 1 4880
box -16 -6 32 210
use FILL  FILL_4190
timestamp 1018054153
transform 1 0 2400 0 1 4880
box -16 -6 32 210
use FILL  FILL_4192
timestamp 1018054153
transform 1 0 2416 0 1 4880
box -16 -6 32 210
use FILL  FILL_4194
timestamp 1018054153
transform 1 0 2432 0 1 4880
box -16 -6 32 210
use FILL  FILL_4196
timestamp 1018054153
transform 1 0 2448 0 1 4880
box -16 -6 32 210
use FILL  FILL_4198
timestamp 1018054153
transform 1 0 2464 0 1 4880
box -16 -6 32 210
use FILL  FILL_4200
timestamp 1018054153
transform 1 0 2480 0 1 4880
box -16 -6 32 210
use FILL  FILL_4202
timestamp 1018054153
transform 1 0 2496 0 1 4880
box -16 -6 32 210
use FILL  FILL_4204
timestamp 1018054153
transform 1 0 2512 0 1 4880
box -16 -6 32 210
use FILL  FILL_4206
timestamp 1018054153
transform 1 0 2528 0 1 4880
box -16 -6 32 210
use FILL  FILL_4208
timestamp 1018054153
transform 1 0 2544 0 1 4880
box -16 -6 32 210
use FILL  FILL_4210
timestamp 1018054153
transform 1 0 2560 0 1 4880
box -16 -6 32 210
use FILL  FILL_4212
timestamp 1018054153
transform 1 0 2576 0 1 4880
box -16 -6 32 210
use FILL  FILL_4214
timestamp 1018054153
transform 1 0 2592 0 1 4880
box -16 -6 32 210
use FILL  FILL_4216
timestamp 1018054153
transform 1 0 2608 0 1 4880
box -16 -6 32 210
use FILL  FILL_4218
timestamp 1018054153
transform 1 0 2624 0 1 4880
box -16 -6 32 210
use FILL  FILL_4220
timestamp 1018054153
transform 1 0 2640 0 1 4880
box -16 -6 32 210
use FILL  FILL_4222
timestamp 1018054153
transform 1 0 2656 0 1 4880
box -16 -6 32 210
use FILL  FILL_4224
timestamp 1018054153
transform 1 0 2672 0 1 4880
box -16 -6 32 210
use FILL  FILL_4226
timestamp 1018054153
transform 1 0 2688 0 1 4880
box -16 -6 32 210
use FILL  FILL_4228
timestamp 1018054153
transform 1 0 2704 0 1 4880
box -16 -6 32 210
use FILL  FILL_4230
timestamp 1018054153
transform 1 0 2720 0 1 4880
box -16 -6 32 210
use FILL  FILL_4232
timestamp 1018054153
transform 1 0 2736 0 1 4880
box -16 -6 32 210
use FILL  FILL_4234
timestamp 1018054153
transform 1 0 2752 0 1 4880
box -16 -6 32 210
use FILL  FILL_4236
timestamp 1018054153
transform 1 0 2768 0 1 4880
box -16 -6 32 210
use FILL  FILL_4238
timestamp 1018054153
transform 1 0 2784 0 1 4880
box -16 -6 32 210
use FILL  FILL_4240
timestamp 1018054153
transform 1 0 2800 0 1 4880
box -16 -6 32 210
use FILL  FILL_4242
timestamp 1018054153
transform 1 0 2816 0 1 4880
box -16 -6 32 210
use FILL  FILL_4244
timestamp 1018054153
transform 1 0 2832 0 1 4880
box -16 -6 32 210
use FILL  FILL_4246
timestamp 1018054153
transform 1 0 2848 0 1 4880
box -16 -6 32 210
use FILL  FILL_4248
timestamp 1018054153
transform 1 0 2864 0 1 4880
box -16 -6 32 210
use FILL  FILL_4250
timestamp 1018054153
transform 1 0 2880 0 1 4880
box -16 -6 32 210
use FILL  FILL_4252
timestamp 1018054153
transform 1 0 2896 0 1 4880
box -16 -6 32 210
use FILL  FILL_4254
timestamp 1018054153
transform 1 0 2912 0 1 4880
box -16 -6 32 210
use FILL  FILL_4256
timestamp 1018054153
transform 1 0 2928 0 1 4880
box -16 -6 32 210
use FILL  FILL_4258
timestamp 1018054153
transform 1 0 2944 0 1 4880
box -16 -6 32 210
use FILL  FILL_4260
timestamp 1018054153
transform 1 0 2960 0 1 4880
box -16 -6 32 210
use FILL  FILL_4262
timestamp 1018054153
transform 1 0 2976 0 1 4880
box -16 -6 32 210
use FILL  FILL_4264
timestamp 1018054153
transform 1 0 2992 0 1 4880
box -16 -6 32 210
use FILL  FILL_4266
timestamp 1018054153
transform 1 0 3008 0 1 4880
box -16 -6 32 210
use FILL  FILL_4268
timestamp 1018054153
transform 1 0 3024 0 1 4880
box -16 -6 32 210
use FILL  FILL_4270
timestamp 1018054153
transform 1 0 3040 0 1 4880
box -16 -6 32 210
use FILL  FILL_4272
timestamp 1018054153
transform 1 0 3056 0 1 4880
box -16 -6 32 210
use FILL  FILL_4274
timestamp 1018054153
transform 1 0 3072 0 1 4880
box -16 -6 32 210
use FILL  FILL_4276
timestamp 1018054153
transform 1 0 3088 0 1 4880
box -16 -6 32 210
use FILL  FILL_4278
timestamp 1018054153
transform 1 0 3104 0 1 4880
box -16 -6 32 210
use FILL  FILL_4280
timestamp 1018054153
transform 1 0 3120 0 1 4880
box -16 -6 32 210
use FILL  FILL_4282
timestamp 1018054153
transform 1 0 3136 0 1 4880
box -16 -6 32 210
use FILL  FILL_4284
timestamp 1018054153
transform 1 0 3152 0 1 4880
box -16 -6 32 210
use FILL  FILL_4286
timestamp 1018054153
transform 1 0 3168 0 1 4880
box -16 -6 32 210
use FILL  FILL_4288
timestamp 1018054153
transform 1 0 3184 0 1 4880
box -16 -6 32 210
use FILL  FILL_4290
timestamp 1018054153
transform 1 0 3200 0 1 4880
box -16 -6 32 210
use FILL  FILL_4292
timestamp 1018054153
transform 1 0 3216 0 1 4880
box -16 -6 32 210
use FILL  FILL_4294
timestamp 1018054153
transform 1 0 3232 0 1 4880
box -16 -6 32 210
use FILL  FILL_4296
timestamp 1018054153
transform 1 0 3248 0 1 4880
box -16 -6 32 210
use FILL  FILL_4298
timestamp 1018054153
transform 1 0 3264 0 1 4880
box -16 -6 32 210
use FILL  FILL_4300
timestamp 1018054153
transform 1 0 3280 0 1 4880
box -16 -6 32 210
use FILL  FILL_4302
timestamp 1018054153
transform 1 0 3296 0 1 4880
box -16 -6 32 210
use FILL  FILL_4304
timestamp 1018054153
transform 1 0 3312 0 1 4880
box -16 -6 32 210
use FILL  FILL_4306
timestamp 1018054153
transform 1 0 3328 0 1 4880
box -16 -6 32 210
use FILL  FILL_4308
timestamp 1018054153
transform 1 0 3344 0 1 4880
box -16 -6 32 210
use FILL  FILL_4310
timestamp 1018054153
transform 1 0 3360 0 1 4880
box -16 -6 32 210
use FILL  FILL_4312
timestamp 1018054153
transform 1 0 3376 0 1 4880
box -16 -6 32 210
use FILL  FILL_4314
timestamp 1018054153
transform 1 0 3392 0 1 4880
box -16 -6 32 210
use FILL  FILL_4316
timestamp 1018054153
transform 1 0 3408 0 1 4880
box -16 -6 32 210
use FILL  FILL_4318
timestamp 1018054153
transform 1 0 3424 0 1 4880
box -16 -6 32 210
use FILL  FILL_4320
timestamp 1018054153
transform 1 0 3440 0 1 4880
box -16 -6 32 210
use FILL  FILL_4322
timestamp 1018054153
transform 1 0 3456 0 1 4880
box -16 -6 32 210
use FILL  FILL_4324
timestamp 1018054153
transform 1 0 3472 0 1 4880
box -16 -6 32 210
use FILL  FILL_4326
timestamp 1018054153
transform 1 0 3488 0 1 4880
box -16 -6 32 210
use FILL  FILL_4328
timestamp 1018054153
transform 1 0 3504 0 1 4880
box -16 -6 32 210
use FILL  FILL_4330
timestamp 1018054153
transform 1 0 3520 0 1 4880
box -16 -6 32 210
use FILL  FILL_4332
timestamp 1018054153
transform 1 0 3536 0 1 4880
box -16 -6 32 210
use FILL  FILL_4334
timestamp 1018054153
transform 1 0 3552 0 1 4880
box -16 -6 32 210
use FILL  FILL_4336
timestamp 1018054153
transform 1 0 3568 0 1 4880
box -16 -6 32 210
use FILL  FILL_4338
timestamp 1018054153
transform 1 0 3584 0 1 4880
box -16 -6 32 210
use FILL  FILL_4340
timestamp 1018054153
transform 1 0 3600 0 1 4880
box -16 -6 32 210
use FILL  FILL_4342
timestamp 1018054153
transform 1 0 3616 0 1 4880
box -16 -6 32 210
use FILL  FILL_4344
timestamp 1018054153
transform 1 0 3632 0 1 4880
box -16 -6 32 210
use FILL  FILL_4346
timestamp 1018054153
transform 1 0 3648 0 1 4880
box -16 -6 32 210
use FILL  FILL_4348
timestamp 1018054153
transform 1 0 3664 0 1 4880
box -16 -6 32 210
use FILL  FILL_4350
timestamp 1018054153
transform 1 0 3680 0 1 4880
box -16 -6 32 210
use FILL  FILL_4352
timestamp 1018054153
transform 1 0 3696 0 1 4880
box -16 -6 32 210
use FILL  FILL_4354
timestamp 1018054153
transform 1 0 3712 0 1 4880
box -16 -6 32 210
use FILL  FILL_4356
timestamp 1018054153
transform 1 0 3728 0 1 4880
box -16 -6 32 210
use FILL  FILL_4358
timestamp 1018054153
transform 1 0 3744 0 1 4880
box -16 -6 32 210
use FILL  FILL_4360
timestamp 1018054153
transform 1 0 3760 0 1 4880
box -16 -6 32 210
use FILL  FILL_4362
timestamp 1018054153
transform 1 0 3776 0 1 4880
box -16 -6 32 210
use INVX2  INVX2_0
timestamp 1053022145
transform 1 0 3792 0 1 4880
box -18 -6 52 210
use FILL  FILL_4364
timestamp 1018054153
transform 1 0 3824 0 1 4880
box -16 -6 32 210
use FILL  FILL_4368
timestamp 1018054153
transform 1 0 3840 0 1 4880
box -16 -6 32 210
use FILL  FILL_4370
timestamp 1018054153
transform 1 0 3856 0 1 4880
box -16 -6 32 210
use FILL  FILL_4372
timestamp 1018054153
transform 1 0 3872 0 1 4880
box -16 -6 32 210
use FILL  FILL_4374
timestamp 1018054153
transform 1 0 3888 0 1 4880
box -16 -6 32 210
use FILL  FILL_4376
timestamp 1018054153
transform 1 0 3904 0 1 4880
box -16 -6 32 210
use FILL  FILL_4378
timestamp 1018054153
transform 1 0 3920 0 1 4880
box -16 -6 32 210
use FILL  FILL_4380
timestamp 1018054153
transform 1 0 3936 0 1 4880
box -16 -6 32 210
use FILL  FILL_4382
timestamp 1018054153
transform 1 0 3952 0 1 4880
box -16 -6 32 210
use FILL  FILL_4384
timestamp 1018054153
transform 1 0 3968 0 1 4880
box -16 -6 32 210
use FILL  FILL_4386
timestamp 1018054153
transform 1 0 3984 0 1 4880
box -16 -6 32 210
use FILL  FILL_4388
timestamp 1018054153
transform 1 0 4000 0 1 4880
box -16 -6 32 210
use FILL  FILL_4390
timestamp 1018054153
transform 1 0 4016 0 1 4880
box -16 -6 32 210
use FILL  FILL_4392
timestamp 1018054153
transform 1 0 4032 0 1 4880
box -16 -6 32 210
use FILL  FILL_4394
timestamp 1018054153
transform 1 0 4048 0 1 4880
box -16 -6 32 210
use FILL  FILL_4396
timestamp 1018054153
transform 1 0 4064 0 1 4880
box -16 -6 32 210
use FILL  FILL_4398
timestamp 1018054153
transform 1 0 4080 0 1 4880
box -16 -6 32 210
use FILL  FILL_4400
timestamp 1018054153
transform 1 0 4096 0 1 4880
box -16 -6 32 210
use FILL  FILL_4402
timestamp 1018054153
transform 1 0 4112 0 1 4880
box -16 -6 32 210
use FILL  FILL_4404
timestamp 1018054153
transform 1 0 4128 0 1 4880
box -16 -6 32 210
use BUFX2  BUFX2_0
timestamp 1090542073
transform 1 0 4144 0 1 4880
box -10 -6 56 210
use FILL  FILL_4406
timestamp 1018054153
transform 1 0 4192 0 1 4880
box -16 -6 32 210
use FILL  FILL_4411
timestamp 1018054153
transform 1 0 4208 0 1 4880
box -16 -6 32 210
use FILL  FILL_4413
timestamp 1018054153
transform 1 0 4224 0 1 4880
box -16 -6 32 210
use FILL  FILL_4415
timestamp 1018054153
transform 1 0 4240 0 1 4880
box -16 -6 32 210
use FILL  FILL_4417
timestamp 1018054153
transform 1 0 4256 0 1 4880
box -16 -6 32 210
use FILL  FILL_4419
timestamp 1018054153
transform 1 0 4272 0 1 4880
box -16 -6 32 210
use FILL  FILL_4421
timestamp 1018054153
transform 1 0 4288 0 1 4880
box -16 -6 32 210
use FILL  FILL_4423
timestamp 1018054153
transform 1 0 4304 0 1 4880
box -16 -6 32 210
use FILL  FILL_4425
timestamp 1018054153
transform 1 0 4320 0 1 4880
box -16 -6 32 210
use FILL  FILL_4427
timestamp 1018054153
transform 1 0 4336 0 1 4880
box -16 -6 32 210
use FILL  FILL_4429
timestamp 1018054153
transform 1 0 4352 0 1 4880
box -16 -6 32 210
use FILL  FILL_4431
timestamp 1018054153
transform 1 0 4368 0 1 4880
box -16 -6 32 210
use FILL  FILL_4433
timestamp 1018054153
transform 1 0 4384 0 1 4880
box -16 -6 32 210
use FILL  FILL_4435
timestamp 1018054153
transform 1 0 4400 0 1 4880
box -16 -6 32 210
use FILL  FILL_4437
timestamp 1018054153
transform 1 0 4416 0 1 4880
box -16 -6 32 210
use FILL  FILL_4439
timestamp 1018054153
transform 1 0 4432 0 1 4880
box -16 -6 32 210
use FILL  FILL_4441
timestamp 1018054153
transform 1 0 4448 0 1 4880
box -16 -6 32 210
use FILL  FILL_4443
timestamp 1018054153
transform 1 0 4464 0 1 4880
box -16 -6 32 210
use BUFX2  BUFX2_1
timestamp 1090542073
transform 1 0 4480 0 1 4880
box -10 -6 56 210
use FILL  FILL_4445
timestamp 1018054153
transform 1 0 4528 0 1 4880
box -16 -6 32 210
use FILL  FILL_4450
timestamp 1018054153
transform 1 0 4544 0 1 4880
box -16 -6 32 210
use FILL  FILL_4452
timestamp 1018054153
transform 1 0 4560 0 1 4880
box -16 -6 32 210
use FILL  FILL_4454
timestamp 1018054153
transform 1 0 4576 0 1 4880
box -16 -6 32 210
use FILL  FILL_4456
timestamp 1018054153
transform 1 0 4592 0 1 4880
box -16 -6 32 210
use mult_pad_VIA2  mult_pad_VIA2_4
timestamp 1542725905
transform 1 0 4625 0 1 4880
box -6 -6 6 6
use M2_M1  M2_M1_211
timestamp 1542725905
transform 1 0 6600 0 1 4970
box -4 -4 4 4
use M2_M1  M2_M1_200
timestamp 1542725905
transform 1 0 6872 0 1 4990
box -4 -4 4 4
use PADOUT  PADOUT_0
timestamp 1084294529
transform 0 1 8000 -1 0 5600
box -12 -6 606 2000
use M3_M2  M3_M2_76
timestamp 1542725905
transform 1 0 8002 0 1 4910
box -6 -6 6 6
use M2_M1  M2_M1_221
timestamp 1542725905
transform 1 0 4440 0 1 4710
box -4 -4 4 4
use M3_M2  M3_M2_77
timestamp 1542725905
transform 1 0 5320 0 1 4870
box -6 -6 6 6
use M3_M2  M3_M2_78
timestamp 1542725905
transform 1 0 5400 0 1 4870
box -6 -6 6 6
use M3_M2  M3_M2_79
timestamp 1542725905
transform 1 0 5848 0 1 4870
box -6 -6 6 6
use M3_M2  M3_M2_80
timestamp 1542725905
transform 1 0 6280 0 1 4870
box -6 -6 6 6
use mult_pad_VIA2  mult_pad_VIA2_5
timestamp 1542725905
transform 1 0 6565 0 1 4880
box -6 -6 6 6
use FILL  FILL_4457
timestamp 1018054153
transform 1 0 6592 0 1 4880
box -16 -6 32 210
use FILL  FILL_4460
timestamp 1018054153
transform 1 0 6608 0 1 4880
box -16 -6 32 210
use FILL  FILL_4462
timestamp 1018054153
transform 1 0 6624 0 1 4880
box -16 -6 32 210
use FILL  FILL_4464
timestamp 1018054153
transform 1 0 6640 0 1 4880
box -16 -6 32 210
use FILL  FILL_4466
timestamp 1018054153
transform 1 0 6656 0 1 4880
box -16 -6 32 210
use FILL  FILL_4468
timestamp 1018054153
transform 1 0 6672 0 1 4880
box -16 -6 32 210
use FILL  FILL_4470
timestamp 1018054153
transform 1 0 6688 0 1 4880
box -16 -6 32 210
use FILL  FILL_4472
timestamp 1018054153
transform 1 0 6704 0 1 4880
box -16 -6 32 210
use FILL  FILL_4474
timestamp 1018054153
transform 1 0 6720 0 1 4880
box -16 -6 32 210
use FILL  FILL_4476
timestamp 1018054153
transform 1 0 6736 0 1 4880
box -16 -6 32 210
use FILL  FILL_4478
timestamp 1018054153
transform 1 0 6752 0 1 4880
box -16 -6 32 210
use FILL  FILL_4480
timestamp 1018054153
transform 1 0 6768 0 1 4880
box -16 -6 32 210
use FILL  FILL_4482
timestamp 1018054153
transform 1 0 6784 0 1 4880
box -16 -6 32 210
use FILL  FILL_4484
timestamp 1018054153
transform 1 0 6800 0 1 4880
box -16 -6 32 210
use FILL  FILL_4486
timestamp 1018054153
transform 1 0 6816 0 1 4880
box -16 -6 32 210
use FILL  FILL_4488
timestamp 1018054153
transform 1 0 6832 0 1 4880
box -16 -6 32 210
use FILL  FILL_4490
timestamp 1018054153
transform 1 0 6848 0 1 4880
box -16 -6 32 210
use FILL  FILL_4492
timestamp 1018054153
transform 1 0 6864 0 1 4880
box -16 -6 32 210
use FILL  FILL_4494
timestamp 1018054153
transform 1 0 6880 0 1 4880
box -16 -6 32 210
use FILL  FILL_4496
timestamp 1018054153
transform 1 0 6896 0 1 4880
box -16 -6 32 210
use FILL  FILL_4498
timestamp 1018054153
transform 1 0 6912 0 1 4880
box -16 -6 32 210
use FILL  FILL_4500
timestamp 1018054153
transform 1 0 6928 0 1 4880
box -16 -6 32 210
use FILL  FILL_4502
timestamp 1018054153
transform 1 0 6944 0 1 4880
box -16 -6 32 210
use FILL  FILL_4504
timestamp 1018054153
transform 1 0 6960 0 1 4880
box -16 -6 32 210
use FILL  FILL_4506
timestamp 1018054153
transform 1 0 6976 0 1 4880
box -16 -6 32 210
use FILL  FILL_4508
timestamp 1018054153
transform 1 0 6992 0 1 4880
box -16 -6 32 210
use FILL  FILL_4510
timestamp 1018054153
transform 1 0 7008 0 1 4880
box -16 -6 32 210
use FILL  FILL_4512
timestamp 1018054153
transform 1 0 7024 0 1 4880
box -16 -6 32 210
use FILL  FILL_4514
timestamp 1018054153
transform 1 0 7040 0 1 4880
box -16 -6 32 210
use FILL  FILL_4516
timestamp 1018054153
transform 1 0 7056 0 1 4880
box -16 -6 32 210
use FILL  FILL_4518
timestamp 1018054153
transform 1 0 7072 0 1 4880
box -16 -6 32 210
use FILL  FILL_4520
timestamp 1018054153
transform 1 0 7088 0 1 4880
box -16 -6 32 210
use FILL  FILL_4522
timestamp 1018054153
transform 1 0 7104 0 1 4880
box -16 -6 32 210
use FILL  FILL_4524
timestamp 1018054153
transform 1 0 7120 0 1 4880
box -16 -6 32 210
use FILL  FILL_4526
timestamp 1018054153
transform 1 0 7136 0 1 4880
box -16 -6 32 210
use FILL  FILL_4528
timestamp 1018054153
transform 1 0 7152 0 1 4880
box -16 -6 32 210
use FILL  FILL_4530
timestamp 1018054153
transform 1 0 7168 0 1 4880
box -16 -6 32 210
use FILL  FILL_4532
timestamp 1018054153
transform 1 0 7184 0 1 4880
box -16 -6 32 210
use FILL  FILL_4534
timestamp 1018054153
transform 1 0 7200 0 1 4880
box -16 -6 32 210
use FILL  FILL_4536
timestamp 1018054153
transform 1 0 7216 0 1 4880
box -16 -6 32 210
use FILL  FILL_4538
timestamp 1018054153
transform 1 0 7232 0 1 4880
box -16 -6 32 210
use FILL  FILL_4540
timestamp 1018054153
transform 1 0 7248 0 1 4880
box -16 -6 32 210
use FILL  FILL_4542
timestamp 1018054153
transform 1 0 7264 0 1 4880
box -16 -6 32 210
use FILL  FILL_4544
timestamp 1018054153
transform 1 0 7280 0 1 4880
box -16 -6 32 210
use FILL  FILL_4546
timestamp 1018054153
transform 1 0 7296 0 1 4880
box -16 -6 32 210
use FILL  FILL_4548
timestamp 1018054153
transform 1 0 7312 0 1 4880
box -16 -6 32 210
use FILL  FILL_4550
timestamp 1018054153
transform 1 0 7328 0 1 4880
box -16 -6 32 210
use FILL  FILL_4552
timestamp 1018054153
transform 1 0 7344 0 1 4880
box -16 -6 32 210
use FILL  FILL_4554
timestamp 1018054153
transform 1 0 7360 0 1 4880
box -16 -6 32 210
use FILL  FILL_4556
timestamp 1018054153
transform 1 0 7376 0 1 4880
box -16 -6 32 210
use FILL  FILL_4558
timestamp 1018054153
transform 1 0 7392 0 1 4880
box -16 -6 32 210
use FILL  FILL_4560
timestamp 1018054153
transform 1 0 7408 0 1 4880
box -16 -6 32 210
use FILL  FILL_4562
timestamp 1018054153
transform 1 0 7424 0 1 4880
box -16 -6 32 210
use FILL  FILL_4564
timestamp 1018054153
transform 1 0 7440 0 1 4880
box -16 -6 32 210
use FILL  FILL_4566
timestamp 1018054153
transform 1 0 7456 0 1 4880
box -16 -6 32 210
use FILL  FILL_4568
timestamp 1018054153
transform 1 0 7472 0 1 4880
box -16 -6 32 210
use FILL  FILL_4570
timestamp 1018054153
transform 1 0 7488 0 1 4880
box -16 -6 32 210
use FILL  FILL_4572
timestamp 1018054153
transform 1 0 7504 0 1 4880
box -16 -6 32 210
use FILL  FILL_4574
timestamp 1018054153
transform 1 0 7520 0 1 4880
box -16 -6 32 210
use FILL  FILL_4576
timestamp 1018054153
transform 1 0 7536 0 1 4880
box -16 -6 32 210
use FILL  FILL_4578
timestamp 1018054153
transform 1 0 7552 0 1 4880
box -16 -6 32 210
use FILL  FILL_4580
timestamp 1018054153
transform 1 0 7568 0 1 4880
box -16 -6 32 210
use FILL  FILL_4582
timestamp 1018054153
transform 1 0 7584 0 1 4880
box -16 -6 32 210
use FILL  FILL_4584
timestamp 1018054153
transform 1 0 7600 0 1 4880
box -16 -6 32 210
use FILL  FILL_4586
timestamp 1018054153
transform 1 0 7616 0 1 4880
box -16 -6 32 210
use FILL  FILL_4588
timestamp 1018054153
transform 1 0 7632 0 1 4880
box -16 -6 32 210
use FILL  FILL_4590
timestamp 1018054153
transform 1 0 7648 0 1 4880
box -16 -6 32 210
use FILL  FILL_4592
timestamp 1018054153
transform 1 0 7664 0 1 4880
box -16 -6 32 210
use FILL  FILL_4594
timestamp 1018054153
transform 1 0 7680 0 1 4880
box -16 -6 32 210
use FILL  FILL_4596
timestamp 1018054153
transform 1 0 7696 0 1 4880
box -16 -6 32 210
use FILL  FILL_4598
timestamp 1018054153
transform 1 0 7712 0 1 4880
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_25
timestamp 1542725905
transform 1 0 7908 0 1 4880
box -48 -6 48 6
use M3_M2  M3_M2_81
timestamp 1542725905
transform 1 0 5768 0 1 4810
box -6 -6 6 6
use M3_M2  M3_M2_82
timestamp 1542725905
transform 1 0 5816 0 1 4810
box -6 -6 6 6
use mult_pad_VIA4  mult_pad_VIA4_2
timestamp 1542725905
transform 1 0 4709 0 1 4713
box -10 -10 10 10
use mult_pad_VIA8  mult_pad_VIA8_2
timestamp 1542725905
transform 1 0 4923 0 1 4707
box -4 -4 4 4
use mult_pad_VIA8  mult_pad_VIA8_3
timestamp 1542725905
transform 1 0 6267 0 1 4707
box -4 -4 4 4
use mult_pad_VIA4  mult_pad_VIA4_3
timestamp 1542725905
transform 1 0 6481 0 1 4713
box -10 -10 10 10
use rca8  rca8_0
timestamp 1542725905
transform 1 0 4699 0 1 4699
box 0 0 1792 258
use mult_pad_VIA1  mult_pad_VIA1_26
timestamp 1542725905
transform 1 0 2212 0 1 4680
box -48 -6 48 6
use FILL  FILL_4175
timestamp 1018054153
transform 1 0 2272 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4177
timestamp 1018054153
transform 1 0 2288 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4179
timestamp 1018054153
transform 1 0 2304 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4181
timestamp 1018054153
transform 1 0 2320 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4183
timestamp 1018054153
transform 1 0 2336 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4185
timestamp 1018054153
transform 1 0 2352 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4187
timestamp 1018054153
transform 1 0 2368 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4189
timestamp 1018054153
transform 1 0 2384 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4191
timestamp 1018054153
transform 1 0 2400 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4193
timestamp 1018054153
transform 1 0 2416 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4195
timestamp 1018054153
transform 1 0 2432 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4197
timestamp 1018054153
transform 1 0 2448 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4199
timestamp 1018054153
transform 1 0 2464 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4201
timestamp 1018054153
transform 1 0 2480 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4203
timestamp 1018054153
transform 1 0 2496 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4205
timestamp 1018054153
transform 1 0 2512 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4207
timestamp 1018054153
transform 1 0 2528 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4209
timestamp 1018054153
transform 1 0 2544 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4211
timestamp 1018054153
transform 1 0 2560 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4213
timestamp 1018054153
transform 1 0 2576 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4215
timestamp 1018054153
transform 1 0 2592 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4217
timestamp 1018054153
transform 1 0 2608 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4219
timestamp 1018054153
transform 1 0 2624 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4221
timestamp 1018054153
transform 1 0 2640 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4223
timestamp 1018054153
transform 1 0 2656 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4225
timestamp 1018054153
transform 1 0 2672 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4227
timestamp 1018054153
transform 1 0 2688 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4229
timestamp 1018054153
transform 1 0 2704 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4231
timestamp 1018054153
transform 1 0 2720 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4233
timestamp 1018054153
transform 1 0 2736 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4235
timestamp 1018054153
transform 1 0 2752 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4237
timestamp 1018054153
transform 1 0 2768 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4239
timestamp 1018054153
transform 1 0 2784 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4241
timestamp 1018054153
transform 1 0 2800 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4243
timestamp 1018054153
transform 1 0 2816 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4245
timestamp 1018054153
transform 1 0 2832 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4247
timestamp 1018054153
transform 1 0 2848 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4249
timestamp 1018054153
transform 1 0 2864 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4251
timestamp 1018054153
transform 1 0 2880 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4253
timestamp 1018054153
transform 1 0 2896 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4255
timestamp 1018054153
transform 1 0 2912 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4257
timestamp 1018054153
transform 1 0 2928 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4259
timestamp 1018054153
transform 1 0 2944 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4261
timestamp 1018054153
transform 1 0 2960 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4263
timestamp 1018054153
transform 1 0 2976 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4265
timestamp 1018054153
transform 1 0 2992 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4267
timestamp 1018054153
transform 1 0 3008 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4269
timestamp 1018054153
transform 1 0 3024 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4271
timestamp 1018054153
transform 1 0 3040 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4273
timestamp 1018054153
transform 1 0 3056 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4275
timestamp 1018054153
transform 1 0 3072 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4277
timestamp 1018054153
transform 1 0 3088 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4279
timestamp 1018054153
transform 1 0 3104 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4281
timestamp 1018054153
transform 1 0 3120 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4283
timestamp 1018054153
transform 1 0 3136 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4285
timestamp 1018054153
transform 1 0 3152 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4287
timestamp 1018054153
transform 1 0 3168 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4289
timestamp 1018054153
transform 1 0 3184 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4291
timestamp 1018054153
transform 1 0 3200 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4293
timestamp 1018054153
transform 1 0 3216 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4295
timestamp 1018054153
transform 1 0 3232 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4297
timestamp 1018054153
transform 1 0 3248 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4299
timestamp 1018054153
transform 1 0 3264 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4301
timestamp 1018054153
transform 1 0 3280 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4303
timestamp 1018054153
transform 1 0 3296 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4305
timestamp 1018054153
transform 1 0 3312 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4307
timestamp 1018054153
transform 1 0 3328 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4309
timestamp 1018054153
transform 1 0 3344 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4311
timestamp 1018054153
transform 1 0 3360 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4313
timestamp 1018054153
transform 1 0 3376 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4315
timestamp 1018054153
transform 1 0 3392 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4317
timestamp 1018054153
transform 1 0 3408 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4319
timestamp 1018054153
transform 1 0 3424 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4321
timestamp 1018054153
transform 1 0 3440 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4323
timestamp 1018054153
transform 1 0 3456 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4325
timestamp 1018054153
transform 1 0 3472 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4327
timestamp 1018054153
transform 1 0 3488 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4329
timestamp 1018054153
transform 1 0 3504 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4331
timestamp 1018054153
transform 1 0 3520 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4333
timestamp 1018054153
transform 1 0 3536 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4335
timestamp 1018054153
transform 1 0 3552 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4337
timestamp 1018054153
transform 1 0 3568 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4339
timestamp 1018054153
transform 1 0 3584 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4341
timestamp 1018054153
transform 1 0 3600 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4343
timestamp 1018054153
transform 1 0 3616 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4345
timestamp 1018054153
transform 1 0 3632 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4347
timestamp 1018054153
transform 1 0 3648 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4349
timestamp 1018054153
transform 1 0 3664 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4351
timestamp 1018054153
transform 1 0 3680 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4353
timestamp 1018054153
transform 1 0 3696 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4355
timestamp 1018054153
transform 1 0 3712 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4357
timestamp 1018054153
transform 1 0 3728 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4359
timestamp 1018054153
transform 1 0 3744 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4361
timestamp 1018054153
transform 1 0 3760 0 -1 4880
box -16 -6 32 210
use M2_M1  M2_M1_227
timestamp 1542725905
transform 1 0 3800 0 1 4680
box -4 -4 4 4
use FILL  FILL_4363
timestamp 1018054153
transform 1 0 3776 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4365
timestamp 1018054153
transform 1 0 3792 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4366
timestamp 1018054153
transform 1 0 3808 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4367
timestamp 1018054153
transform 1 0 3824 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4369
timestamp 1018054153
transform 1 0 3840 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4371
timestamp 1018054153
transform 1 0 3856 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4373
timestamp 1018054153
transform 1 0 3872 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4375
timestamp 1018054153
transform 1 0 3888 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4377
timestamp 1018054153
transform 1 0 3904 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4379
timestamp 1018054153
transform 1 0 3920 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4381
timestamp 1018054153
transform 1 0 3936 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4383
timestamp 1018054153
transform 1 0 3952 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4385
timestamp 1018054153
transform 1 0 3968 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4387
timestamp 1018054153
transform 1 0 3984 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4389
timestamp 1018054153
transform 1 0 4000 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4391
timestamp 1018054153
transform 1 0 4016 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4393
timestamp 1018054153
transform 1 0 4032 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4395
timestamp 1018054153
transform 1 0 4048 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4397
timestamp 1018054153
transform 1 0 4064 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4399
timestamp 1018054153
transform 1 0 4080 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4401
timestamp 1018054153
transform 1 0 4096 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4403
timestamp 1018054153
transform 1 0 4112 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4405
timestamp 1018054153
transform 1 0 4128 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4407
timestamp 1018054153
transform 1 0 4144 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4408
timestamp 1018054153
transform 1 0 4160 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4409
timestamp 1018054153
transform 1 0 4176 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4410
timestamp 1018054153
transform 1 0 4192 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4412
timestamp 1018054153
transform 1 0 4208 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4414
timestamp 1018054153
transform 1 0 4224 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4416
timestamp 1018054153
transform 1 0 4240 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4418
timestamp 1018054153
transform 1 0 4256 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4420
timestamp 1018054153
transform 1 0 4272 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4422
timestamp 1018054153
transform 1 0 4288 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4424
timestamp 1018054153
transform 1 0 4304 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4426
timestamp 1018054153
transform 1 0 4320 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4428
timestamp 1018054153
transform 1 0 4336 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4430
timestamp 1018054153
transform 1 0 4352 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4432
timestamp 1018054153
transform 1 0 4368 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4434
timestamp 1018054153
transform 1 0 4384 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4436
timestamp 1018054153
transform 1 0 4400 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4438
timestamp 1018054153
transform 1 0 4416 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4440
timestamp 1018054153
transform 1 0 4432 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4442
timestamp 1018054153
transform 1 0 4448 0 -1 4880
box -16 -6 32 210
use M3_M2  M3_M2_83
timestamp 1542725905
transform 1 0 4488 0 1 4690
box -6 -6 6 6
use FILL  FILL_4444
timestamp 1018054153
transform 1 0 4464 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4446
timestamp 1018054153
transform 1 0 4480 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4447
timestamp 1018054153
transform 1 0 4496 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4448
timestamp 1018054153
transform 1 0 4512 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4449
timestamp 1018054153
transform 1 0 4528 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4451
timestamp 1018054153
transform 1 0 4544 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4453
timestamp 1018054153
transform 1 0 4560 0 -1 4880
box -16 -6 32 210
use M3_M2  M3_M2_84
timestamp 1542725905
transform 1 0 4600 0 1 4690
box -6 -6 6 6
use FILL  FILL_4455
timestamp 1018054153
transform 1 0 4576 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4458
timestamp 1018054153
transform 1 0 4592 0 -1 4880
box -16 -6 32 210
use M2_M1  M2_M1_222
timestamp 1542725905
transform 1 0 4840 0 1 4690
box -4 -4 4 4
use M2_M1  M2_M1_223
timestamp 1542725905
transform 1 0 5224 0 1 4690
box -4 -4 4 4
use M2_M1  M2_M1_224
timestamp 1542725905
transform 1 0 5992 0 1 4690
box -4 -4 4 4
use M2_M1  M2_M1_225
timestamp 1542725905
transform 1 0 6120 0 1 4690
box -4 -4 4 4
use M2_M1  M2_M1_226
timestamp 1542725905
transform 1 0 6520 0 1 4690
box -4 -4 4 4
use mult_pad_VIA2  mult_pad_VIA2_6
timestamp 1542725905
transform 1 0 4649 0 1 4680
box -6 -6 6 6
use mult_pad_VIA2  mult_pad_VIA2_7
timestamp 1542725905
transform 1 0 6541 0 1 4680
box -6 -6 6 6
use M3_M2  M3_M2_85
timestamp 1542725905
transform 1 0 3944 0 1 4630
box -6 -6 6 6
use M2_M1  M2_M1_231
timestamp 1542725905
transform 1 0 4120 0 1 4610
box -4 -4 4 4
use M2_M1  M2_M1_232
timestamp 1542725905
transform 1 0 3800 0 1 4590
box -4 -4 4 4
use M2_M1  M2_M1_233
timestamp 1542725905
transform 1 0 3848 0 1 4570
box -4 -4 4 4
use M2_M1  M2_M1_234
timestamp 1542725905
transform 1 0 3912 0 1 4550
box -4 -4 4 4
use M3_M2  M3_M2_87
timestamp 1542725905
transform 1 0 3912 0 1 4530
box -6 -6 6 6
use M2_M1  M2_M1_235
timestamp 1542725905
transform 1 0 3944 0 1 4530
box -4 -4 4 4
use M3_M2  M3_M2_86
timestamp 1542725905
transform 1 0 4152 0 1 4630
box -6 -6 6 6
use M2_M1  M2_M1_228
timestamp 1542725905
transform 1 0 5144 0 1 4670
box -4 -4 4 4
use M2_M1  M2_M1_229
timestamp 1542725905
transform 1 0 5528 0 1 4670
box -4 -4 4 4
use M2_M1  M2_M1_230
timestamp 1542725905
transform 1 0 6408 0 1 4670
box -4 -4 4 4
use FILL  FILL_4459
timestamp 1018054153
transform 1 0 6592 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4461
timestamp 1018054153
transform 1 0 6608 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4463
timestamp 1018054153
transform 1 0 6624 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4465
timestamp 1018054153
transform 1 0 6640 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4467
timestamp 1018054153
transform 1 0 6656 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4469
timestamp 1018054153
transform 1 0 6672 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4471
timestamp 1018054153
transform 1 0 6688 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4473
timestamp 1018054153
transform 1 0 6704 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4475
timestamp 1018054153
transform 1 0 6720 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4477
timestamp 1018054153
transform 1 0 6736 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4479
timestamp 1018054153
transform 1 0 6752 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4481
timestamp 1018054153
transform 1 0 6768 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4483
timestamp 1018054153
transform 1 0 6784 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4485
timestamp 1018054153
transform 1 0 6800 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4487
timestamp 1018054153
transform 1 0 6816 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4489
timestamp 1018054153
transform 1 0 6832 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4491
timestamp 1018054153
transform 1 0 6848 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4493
timestamp 1018054153
transform 1 0 6864 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4495
timestamp 1018054153
transform 1 0 6880 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4497
timestamp 1018054153
transform 1 0 6896 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4499
timestamp 1018054153
transform 1 0 6912 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4501
timestamp 1018054153
transform 1 0 6928 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4503
timestamp 1018054153
transform 1 0 6944 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4505
timestamp 1018054153
transform 1 0 6960 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4507
timestamp 1018054153
transform 1 0 6976 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4509
timestamp 1018054153
transform 1 0 6992 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4511
timestamp 1018054153
transform 1 0 7008 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4513
timestamp 1018054153
transform 1 0 7024 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4515
timestamp 1018054153
transform 1 0 7040 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4517
timestamp 1018054153
transform 1 0 7056 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4519
timestamp 1018054153
transform 1 0 7072 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4521
timestamp 1018054153
transform 1 0 7088 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4523
timestamp 1018054153
transform 1 0 7104 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4525
timestamp 1018054153
transform 1 0 7120 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4527
timestamp 1018054153
transform 1 0 7136 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4529
timestamp 1018054153
transform 1 0 7152 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4531
timestamp 1018054153
transform 1 0 7168 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4533
timestamp 1018054153
transform 1 0 7184 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4535
timestamp 1018054153
transform 1 0 7200 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4537
timestamp 1018054153
transform 1 0 7216 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4539
timestamp 1018054153
transform 1 0 7232 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4541
timestamp 1018054153
transform 1 0 7248 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4543
timestamp 1018054153
transform 1 0 7264 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4545
timestamp 1018054153
transform 1 0 7280 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4547
timestamp 1018054153
transform 1 0 7296 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4549
timestamp 1018054153
transform 1 0 7312 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4551
timestamp 1018054153
transform 1 0 7328 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4553
timestamp 1018054153
transform 1 0 7344 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4555
timestamp 1018054153
transform 1 0 7360 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4557
timestamp 1018054153
transform 1 0 7376 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4559
timestamp 1018054153
transform 1 0 7392 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4561
timestamp 1018054153
transform 1 0 7408 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4563
timestamp 1018054153
transform 1 0 7424 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4565
timestamp 1018054153
transform 1 0 7440 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4567
timestamp 1018054153
transform 1 0 7456 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4569
timestamp 1018054153
transform 1 0 7472 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4571
timestamp 1018054153
transform 1 0 7488 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4573
timestamp 1018054153
transform 1 0 7504 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4575
timestamp 1018054153
transform 1 0 7520 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4577
timestamp 1018054153
transform 1 0 7536 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4579
timestamp 1018054153
transform 1 0 7552 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4581
timestamp 1018054153
transform 1 0 7568 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4583
timestamp 1018054153
transform 1 0 7584 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4585
timestamp 1018054153
transform 1 0 7600 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4587
timestamp 1018054153
transform 1 0 7616 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4589
timestamp 1018054153
transform 1 0 7632 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4591
timestamp 1018054153
transform 1 0 7648 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4593
timestamp 1018054153
transform 1 0 7664 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4595
timestamp 1018054153
transform 1 0 7680 0 -1 4880
box -16 -6 32 210
use FILL  FILL_4597
timestamp 1018054153
transform 1 0 7696 0 -1 4880
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_27
timestamp 1542725905
transform 1 0 7788 0 1 4680
box -48 -6 48 6
use FILL  FILL_4599
timestamp 1018054153
transform 1 0 7712 0 -1 4880
box -16 -6 32 210
use mult_pad_VIA2  mult_pad_VIA2_8
timestamp 1542725905
transform 1 0 4649 0 1 4649
box -6 -6 6 6
use mult_pad_VIA10  mult_pad_VIA10_0
timestamp 1542725905
transform 1 0 4923 0 1 4649
box -4 -6 4 6
use mult_pad_VIA10  mult_pad_VIA10_1
timestamp 1542725905
transform 1 0 6267 0 1 4649
box -4 -6 4 6
use mult_pad_VIA2  mult_pad_VIA2_9
timestamp 1542725905
transform 1 0 6541 0 1 4649
box -6 -6 6 6
use mult_pad_VIA2  mult_pad_VIA2_10
timestamp 1542725905
transform 1 0 4625 0 1 4625
box -6 -6 6 6
use mult_pad_VIA3  mult_pad_VIA3_2
timestamp 1542725905
transform 1 0 4709 0 1 4625
box -10 -6 10 6
use mult_pad_VIA3  mult_pad_VIA3_3
timestamp 1542725905
transform 1 0 6481 0 1 4625
box -10 -6 10 6
use mult_pad_VIA2  mult_pad_VIA2_11
timestamp 1542725905
transform 1 0 6565 0 1 4625
box -6 -6 6 6
use M3_M2  M3_M2_88
timestamp 1542725905
transform 1 0 4840 0 1 4530
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_28
timestamp 1542725905
transform 1 0 2092 0 1 4480
box -48 -6 48 6
use FILL  FILL_4600
timestamp 1018054153
transform 1 0 2272 0 1 4480
box -16 -6 32 210
use FILL  FILL_4602
timestamp 1018054153
transform 1 0 2288 0 1 4480
box -16 -6 32 210
use FILL  FILL_4604
timestamp 1018054153
transform 1 0 2304 0 1 4480
box -16 -6 32 210
use FILL  FILL_4606
timestamp 1018054153
transform 1 0 2320 0 1 4480
box -16 -6 32 210
use FILL  FILL_4608
timestamp 1018054153
transform 1 0 2336 0 1 4480
box -16 -6 32 210
use FILL  FILL_4610
timestamp 1018054153
transform 1 0 2352 0 1 4480
box -16 -6 32 210
use FILL  FILL_4612
timestamp 1018054153
transform 1 0 2368 0 1 4480
box -16 -6 32 210
use FILL  FILL_4614
timestamp 1018054153
transform 1 0 2384 0 1 4480
box -16 -6 32 210
use FILL  FILL_4616
timestamp 1018054153
transform 1 0 2400 0 1 4480
box -16 -6 32 210
use FILL  FILL_4618
timestamp 1018054153
transform 1 0 2416 0 1 4480
box -16 -6 32 210
use FILL  FILL_4620
timestamp 1018054153
transform 1 0 2432 0 1 4480
box -16 -6 32 210
use FILL  FILL_4622
timestamp 1018054153
transform 1 0 2448 0 1 4480
box -16 -6 32 210
use FILL  FILL_4624
timestamp 1018054153
transform 1 0 2464 0 1 4480
box -16 -6 32 210
use FILL  FILL_4626
timestamp 1018054153
transform 1 0 2480 0 1 4480
box -16 -6 32 210
use FILL  FILL_4628
timestamp 1018054153
transform 1 0 2496 0 1 4480
box -16 -6 32 210
use FILL  FILL_4630
timestamp 1018054153
transform 1 0 2512 0 1 4480
box -16 -6 32 210
use FILL  FILL_4632
timestamp 1018054153
transform 1 0 2528 0 1 4480
box -16 -6 32 210
use FILL  FILL_4634
timestamp 1018054153
transform 1 0 2544 0 1 4480
box -16 -6 32 210
use FILL  FILL_4636
timestamp 1018054153
transform 1 0 2560 0 1 4480
box -16 -6 32 210
use FILL  FILL_4638
timestamp 1018054153
transform 1 0 2576 0 1 4480
box -16 -6 32 210
use FILL  FILL_4640
timestamp 1018054153
transform 1 0 2592 0 1 4480
box -16 -6 32 210
use FILL  FILL_4642
timestamp 1018054153
transform 1 0 2608 0 1 4480
box -16 -6 32 210
use FILL  FILL_4644
timestamp 1018054153
transform 1 0 2624 0 1 4480
box -16 -6 32 210
use FILL  FILL_4646
timestamp 1018054153
transform 1 0 2640 0 1 4480
box -16 -6 32 210
use FILL  FILL_4648
timestamp 1018054153
transform 1 0 2656 0 1 4480
box -16 -6 32 210
use FILL  FILL_4650
timestamp 1018054153
transform 1 0 2672 0 1 4480
box -16 -6 32 210
use FILL  FILL_4652
timestamp 1018054153
transform 1 0 2688 0 1 4480
box -16 -6 32 210
use FILL  FILL_4654
timestamp 1018054153
transform 1 0 2704 0 1 4480
box -16 -6 32 210
use FILL  FILL_4656
timestamp 1018054153
transform 1 0 2720 0 1 4480
box -16 -6 32 210
use FILL  FILL_4658
timestamp 1018054153
transform 1 0 2736 0 1 4480
box -16 -6 32 210
use FILL  FILL_4660
timestamp 1018054153
transform 1 0 2752 0 1 4480
box -16 -6 32 210
use FILL  FILL_4662
timestamp 1018054153
transform 1 0 2768 0 1 4480
box -16 -6 32 210
use FILL  FILL_4664
timestamp 1018054153
transform 1 0 2784 0 1 4480
box -16 -6 32 210
use FILL  FILL_4666
timestamp 1018054153
transform 1 0 2800 0 1 4480
box -16 -6 32 210
use FILL  FILL_4668
timestamp 1018054153
transform 1 0 2816 0 1 4480
box -16 -6 32 210
use FILL  FILL_4670
timestamp 1018054153
transform 1 0 2832 0 1 4480
box -16 -6 32 210
use FILL  FILL_4672
timestamp 1018054153
transform 1 0 2848 0 1 4480
box -16 -6 32 210
use FILL  FILL_4674
timestamp 1018054153
transform 1 0 2864 0 1 4480
box -16 -6 32 210
use FILL  FILL_4676
timestamp 1018054153
transform 1 0 2880 0 1 4480
box -16 -6 32 210
use FILL  FILL_4678
timestamp 1018054153
transform 1 0 2896 0 1 4480
box -16 -6 32 210
use FILL  FILL_4680
timestamp 1018054153
transform 1 0 2912 0 1 4480
box -16 -6 32 210
use FILL  FILL_4682
timestamp 1018054153
transform 1 0 2928 0 1 4480
box -16 -6 32 210
use FILL  FILL_4684
timestamp 1018054153
transform 1 0 2944 0 1 4480
box -16 -6 32 210
use FILL  FILL_4686
timestamp 1018054153
transform 1 0 2960 0 1 4480
box -16 -6 32 210
use FILL  FILL_4688
timestamp 1018054153
transform 1 0 2976 0 1 4480
box -16 -6 32 210
use FILL  FILL_4690
timestamp 1018054153
transform 1 0 2992 0 1 4480
box -16 -6 32 210
use FILL  FILL_4692
timestamp 1018054153
transform 1 0 3008 0 1 4480
box -16 -6 32 210
use FILL  FILL_4694
timestamp 1018054153
transform 1 0 3024 0 1 4480
box -16 -6 32 210
use FILL  FILL_4696
timestamp 1018054153
transform 1 0 3040 0 1 4480
box -16 -6 32 210
use FILL  FILL_4698
timestamp 1018054153
transform 1 0 3056 0 1 4480
box -16 -6 32 210
use FILL  FILL_4700
timestamp 1018054153
transform 1 0 3072 0 1 4480
box -16 -6 32 210
use FILL  FILL_4702
timestamp 1018054153
transform 1 0 3088 0 1 4480
box -16 -6 32 210
use FILL  FILL_4704
timestamp 1018054153
transform 1 0 3104 0 1 4480
box -16 -6 32 210
use FILL  FILL_4706
timestamp 1018054153
transform 1 0 3120 0 1 4480
box -16 -6 32 210
use FILL  FILL_4708
timestamp 1018054153
transform 1 0 3136 0 1 4480
box -16 -6 32 210
use FILL  FILL_4710
timestamp 1018054153
transform 1 0 3152 0 1 4480
box -16 -6 32 210
use FILL  FILL_4712
timestamp 1018054153
transform 1 0 3168 0 1 4480
box -16 -6 32 210
use FILL  FILL_4714
timestamp 1018054153
transform 1 0 3184 0 1 4480
box -16 -6 32 210
use FILL  FILL_4716
timestamp 1018054153
transform 1 0 3200 0 1 4480
box -16 -6 32 210
use FILL  FILL_4718
timestamp 1018054153
transform 1 0 3216 0 1 4480
box -16 -6 32 210
use FILL  FILL_4720
timestamp 1018054153
transform 1 0 3232 0 1 4480
box -16 -6 32 210
use FILL  FILL_4722
timestamp 1018054153
transform 1 0 3248 0 1 4480
box -16 -6 32 210
use FILL  FILL_4724
timestamp 1018054153
transform 1 0 3264 0 1 4480
box -16 -6 32 210
use FILL  FILL_4726
timestamp 1018054153
transform 1 0 3280 0 1 4480
box -16 -6 32 210
use FILL  FILL_4728
timestamp 1018054153
transform 1 0 3296 0 1 4480
box -16 -6 32 210
use FILL  FILL_4730
timestamp 1018054153
transform 1 0 3312 0 1 4480
box -16 -6 32 210
use FILL  FILL_4732
timestamp 1018054153
transform 1 0 3328 0 1 4480
box -16 -6 32 210
use FILL  FILL_4734
timestamp 1018054153
transform 1 0 3344 0 1 4480
box -16 -6 32 210
use FILL  FILL_4736
timestamp 1018054153
transform 1 0 3360 0 1 4480
box -16 -6 32 210
use FILL  FILL_4738
timestamp 1018054153
transform 1 0 3376 0 1 4480
box -16 -6 32 210
use FILL  FILL_4740
timestamp 1018054153
transform 1 0 3392 0 1 4480
box -16 -6 32 210
use FILL  FILL_4742
timestamp 1018054153
transform 1 0 3408 0 1 4480
box -16 -6 32 210
use FILL  FILL_4744
timestamp 1018054153
transform 1 0 3424 0 1 4480
box -16 -6 32 210
use FILL  FILL_4746
timestamp 1018054153
transform 1 0 3440 0 1 4480
box -16 -6 32 210
use FILL  FILL_4748
timestamp 1018054153
transform 1 0 3456 0 1 4480
box -16 -6 32 210
use FILL  FILL_4750
timestamp 1018054153
transform 1 0 3472 0 1 4480
box -16 -6 32 210
use FILL  FILL_4752
timestamp 1018054153
transform 1 0 3488 0 1 4480
box -16 -6 32 210
use FILL  FILL_4754
timestamp 1018054153
transform 1 0 3504 0 1 4480
box -16 -6 32 210
use FILL  FILL_4756
timestamp 1018054153
transform 1 0 3520 0 1 4480
box -16 -6 32 210
use FILL  FILL_4758
timestamp 1018054153
transform 1 0 3536 0 1 4480
box -16 -6 32 210
use FILL  FILL_4760
timestamp 1018054153
transform 1 0 3552 0 1 4480
box -16 -6 32 210
use FILL  FILL_4762
timestamp 1018054153
transform 1 0 3568 0 1 4480
box -16 -6 32 210
use FILL  FILL_4764
timestamp 1018054153
transform 1 0 3584 0 1 4480
box -16 -6 32 210
use FILL  FILL_4766
timestamp 1018054153
transform 1 0 3600 0 1 4480
box -16 -6 32 210
use FILL  FILL_4768
timestamp 1018054153
transform 1 0 3616 0 1 4480
box -16 -6 32 210
use FILL  FILL_4770
timestamp 1018054153
transform 1 0 3632 0 1 4480
box -16 -6 32 210
use FILL  FILL_4772
timestamp 1018054153
transform 1 0 3648 0 1 4480
box -16 -6 32 210
use FILL  FILL_4774
timestamp 1018054153
transform 1 0 3664 0 1 4480
box -16 -6 32 210
use FILL  FILL_4776
timestamp 1018054153
transform 1 0 3680 0 1 4480
box -16 -6 32 210
use FILL  FILL_4778
timestamp 1018054153
transform 1 0 3696 0 1 4480
box -16 -6 32 210
use FILL  FILL_4780
timestamp 1018054153
transform 1 0 3712 0 1 4480
box -16 -6 32 210
use FILL  FILL_4782
timestamp 1018054153
transform 1 0 3728 0 1 4480
box -16 -6 32 210
use FILL  FILL_4784
timestamp 1018054153
transform 1 0 3744 0 1 4480
box -16 -6 32 210
use FILL  FILL_4786
timestamp 1018054153
transform 1 0 3760 0 1 4480
box -16 -6 32 210
use DFFSR  DFFSR_0
timestamp 1071163401
transform 1 0 3776 0 1 4480
box -16 -6 368 210
use FILL  FILL_4788
timestamp 1018054153
transform 1 0 4128 0 1 4480
box -16 -6 32 210
use FILL  FILL_4812
timestamp 1018054153
transform 1 0 4144 0 1 4480
box -16 -6 32 210
use FILL  FILL_4814
timestamp 1018054153
transform 1 0 4160 0 1 4480
box -16 -6 32 210
use FILL  FILL_4816
timestamp 1018054153
transform 1 0 4176 0 1 4480
box -16 -6 32 210
use FILL  FILL_4818
timestamp 1018054153
transform 1 0 4192 0 1 4480
box -16 -6 32 210
use FILL  FILL_4820
timestamp 1018054153
transform 1 0 4208 0 1 4480
box -16 -6 32 210
use FILL  FILL_4822
timestamp 1018054153
transform 1 0 4224 0 1 4480
box -16 -6 32 210
use FILL  FILL_4824
timestamp 1018054153
transform 1 0 4240 0 1 4480
box -16 -6 32 210
use FILL  FILL_4826
timestamp 1018054153
transform 1 0 4256 0 1 4480
box -16 -6 32 210
use FILL  FILL_4828
timestamp 1018054153
transform 1 0 4272 0 1 4480
box -16 -6 32 210
use FILL  FILL_4829
timestamp 1018054153
transform 1 0 4288 0 1 4480
box -16 -6 32 210
use FILL  FILL_4830
timestamp 1018054153
transform 1 0 4304 0 1 4480
box -16 -6 32 210
use FILL  FILL_4831
timestamp 1018054153
transform 1 0 4320 0 1 4480
box -16 -6 32 210
use FILL  FILL_4832
timestamp 1018054153
transform 1 0 4336 0 1 4480
box -16 -6 32 210
use FILL  FILL_4833
timestamp 1018054153
transform 1 0 4352 0 1 4480
box -16 -6 32 210
use FILL  FILL_4834
timestamp 1018054153
transform 1 0 4368 0 1 4480
box -16 -6 32 210
use FILL  FILL_4835
timestamp 1018054153
transform 1 0 4384 0 1 4480
box -16 -6 32 210
use FILL  FILL_4836
timestamp 1018054153
transform 1 0 4400 0 1 4480
box -16 -6 32 210
use FILL  FILL_4837
timestamp 1018054153
transform 1 0 4416 0 1 4480
box -16 -6 32 210
use FILL  FILL_4838
timestamp 1018054153
transform 1 0 4432 0 1 4480
box -16 -6 32 210
use FILL  FILL_4839
timestamp 1018054153
transform 1 0 4448 0 1 4480
box -16 -6 32 210
use FILL  FILL_4840
timestamp 1018054153
transform 1 0 4464 0 1 4480
box -16 -6 32 210
use FILL  FILL_4841
timestamp 1018054153
transform 1 0 4480 0 1 4480
box -16 -6 32 210
use FILL  FILL_4842
timestamp 1018054153
transform 1 0 4496 0 1 4480
box -16 -6 32 210
use FILL  FILL_4843
timestamp 1018054153
transform 1 0 4512 0 1 4480
box -16 -6 32 210
use FILL  FILL_4844
timestamp 1018054153
transform 1 0 4528 0 1 4480
box -16 -6 32 210
use FILL  FILL_4845
timestamp 1018054153
transform 1 0 4544 0 1 4480
box -16 -6 32 210
use FILL  FILL_4846
timestamp 1018054153
transform 1 0 4560 0 1 4480
box -16 -6 32 210
use FILL  FILL_4847
timestamp 1018054153
transform 1 0 4576 0 1 4480
box -16 -6 32 210
use FILL  FILL_4848
timestamp 1018054153
transform 1 0 4592 0 1 4480
box -16 -6 32 210
use PADINC  PADINC_7
timestamp 1084294328
transform 0 -1 2000 1 0 4400
box -12 -6 606 2000
use M3_M2  M3_M2_92
timestamp 1542725905
transform 1 0 1998 0 1 4330
box -6 -6 6 6
use M3_M2  M3_M2_93
timestamp 1542725905
transform 1 0 3048 0 1 4330
box -6 -6 6 6
use M3_M2  M3_M2_89
timestamp 1542725905
transform 1 0 3848 0 1 4410
box -6 -6 6 6
use M2_M1  M2_M1_236
timestamp 1542725905
transform 1 0 4440 0 1 4430
box -4 -4 4 4
use M3_M2  M3_M2_90
timestamp 1542725905
transform 1 0 4344 0 1 4410
box -6 -6 6 6
use M2_M1  M2_M1_239
timestamp 1542725905
transform 1 0 4408 0 1 4410
box -4 -4 4 4
use M2_M1  M2_M1_244
timestamp 1542725905
transform 1 0 4344 0 1 4390
box -4 -4 4 4
use M2_M1  M2_M1_247
timestamp 1542725905
transform 1 0 4296 0 1 4370
box -4 -4 4 4
use M2_M1  M2_M1_250
timestamp 1542725905
transform 1 0 4600 0 1 4350
box -4 -4 4 4
use M2_M1  M2_M1_237
timestamp 1542725905
transform 1 0 5256 0 1 4430
box -4 -4 4 4
use M3_M2  M3_M2_91
timestamp 1542725905
transform 1 0 5096 0 1 4410
box -6 -6 6 6
use M2_M1  M2_M1_240
timestamp 1542725905
transform 1 0 5224 0 1 4410
box -4 -4 4 4
use M2_M1  M2_M1_245
timestamp 1542725905
transform 1 0 5160 0 1 4390
box -4 -4 4 4
use M2_M1  M2_M1_248
timestamp 1542725905
transform 1 0 5128 0 1 4370
box -4 -4 4 4
use M2_M1  M2_M1_251
timestamp 1542725905
transform 1 0 5416 0 1 4350
box -4 -4 4 4
use M3_M2  M3_M2_94
timestamp 1542725905
transform 1 0 5112 0 1 4310
box -6 -6 6 6
use M3_M2  M3_M2_95
timestamp 1542725905
transform 1 0 5160 0 1 4310
box -6 -6 6 6
use M3_M2  M3_M2_96
timestamp 1542725905
transform 1 0 5416 0 1 4310
box -6 -6 6 6
use M2_M1  M2_M1_238
timestamp 1542725905
transform 1 0 6168 0 1 4430
box -4 -4 4 4
use M2_M1  M2_M1_241
timestamp 1542725905
transform 1 0 6136 0 1 4410
box -4 -4 4 4
use M2_M1  M2_M1_246
timestamp 1542725905
transform 1 0 6072 0 1 4390
box -4 -4 4 4
use M2_M1  M2_M1_249
timestamp 1542725905
transform 1 0 6040 0 1 4370
box -4 -4 4 4
use FILL  FILL_4849
timestamp 1018054153
transform 1 0 6592 0 1 4480
box -16 -6 32 210
use FILL  FILL_4930
timestamp 1018054153
transform 1 0 6608 0 1 4480
box -16 -6 32 210
use FILL  FILL_4932
timestamp 1018054153
transform 1 0 6624 0 1 4480
box -16 -6 32 210
use FILL  FILL_4934
timestamp 1018054153
transform 1 0 6640 0 1 4480
box -16 -6 32 210
use FILL  FILL_4936
timestamp 1018054153
transform 1 0 6656 0 1 4480
box -16 -6 32 210
use FILL  FILL_4938
timestamp 1018054153
transform 1 0 6672 0 1 4480
box -16 -6 32 210
use FILL  FILL_4940
timestamp 1018054153
transform 1 0 6688 0 1 4480
box -16 -6 32 210
use FILL  FILL_4942
timestamp 1018054153
transform 1 0 6704 0 1 4480
box -16 -6 32 210
use FILL  FILL_4944
timestamp 1018054153
transform 1 0 6720 0 1 4480
box -16 -6 32 210
use FILL  FILL_4946
timestamp 1018054153
transform 1 0 6736 0 1 4480
box -16 -6 32 210
use FILL  FILL_4948
timestamp 1018054153
transform 1 0 6752 0 1 4480
box -16 -6 32 210
use FILL  FILL_4950
timestamp 1018054153
transform 1 0 6768 0 1 4480
box -16 -6 32 210
use FILL  FILL_4952
timestamp 1018054153
transform 1 0 6784 0 1 4480
box -16 -6 32 210
use FILL  FILL_4954
timestamp 1018054153
transform 1 0 6800 0 1 4480
box -16 -6 32 210
use FILL  FILL_4956
timestamp 1018054153
transform 1 0 6816 0 1 4480
box -16 -6 32 210
use FILL  FILL_4958
timestamp 1018054153
transform 1 0 6832 0 1 4480
box -16 -6 32 210
use FILL  FILL_4959
timestamp 1018054153
transform 1 0 6848 0 1 4480
box -16 -6 32 210
use FILL  FILL_4960
timestamp 1018054153
transform 1 0 6864 0 1 4480
box -16 -6 32 210
use FILL  FILL_4961
timestamp 1018054153
transform 1 0 6880 0 1 4480
box -16 -6 32 210
use FILL  FILL_4963
timestamp 1018054153
transform 1 0 6896 0 1 4480
box -16 -6 32 210
use FILL  FILL_4965
timestamp 1018054153
transform 1 0 6912 0 1 4480
box -16 -6 32 210
use FILL  FILL_4967
timestamp 1018054153
transform 1 0 6928 0 1 4480
box -16 -6 32 210
use FILL  FILL_4969
timestamp 1018054153
transform 1 0 6944 0 1 4480
box -16 -6 32 210
use FILL  FILL_4971
timestamp 1018054153
transform 1 0 6960 0 1 4480
box -16 -6 32 210
use FILL  FILL_4973
timestamp 1018054153
transform 1 0 6976 0 1 4480
box -16 -6 32 210
use FILL  FILL_4975
timestamp 1018054153
transform 1 0 6992 0 1 4480
box -16 -6 32 210
use FILL  FILL_4977
timestamp 1018054153
transform 1 0 7008 0 1 4480
box -16 -6 32 210
use FILL  FILL_4979
timestamp 1018054153
transform 1 0 7024 0 1 4480
box -16 -6 32 210
use FILL  FILL_4981
timestamp 1018054153
transform 1 0 7040 0 1 4480
box -16 -6 32 210
use FILL  FILL_4983
timestamp 1018054153
transform 1 0 7056 0 1 4480
box -16 -6 32 210
use FILL  FILL_4985
timestamp 1018054153
transform 1 0 7072 0 1 4480
box -16 -6 32 210
use FILL  FILL_4987
timestamp 1018054153
transform 1 0 7088 0 1 4480
box -16 -6 32 210
use FILL  FILL_4989
timestamp 1018054153
transform 1 0 7104 0 1 4480
box -16 -6 32 210
use FILL  FILL_4991
timestamp 1018054153
transform 1 0 7120 0 1 4480
box -16 -6 32 210
use FILL  FILL_4993
timestamp 1018054153
transform 1 0 7136 0 1 4480
box -16 -6 32 210
use FILL  FILL_4995
timestamp 1018054153
transform 1 0 7152 0 1 4480
box -16 -6 32 210
use FILL  FILL_4997
timestamp 1018054153
transform 1 0 7168 0 1 4480
box -16 -6 32 210
use FILL  FILL_4999
timestamp 1018054153
transform 1 0 7184 0 1 4480
box -16 -6 32 210
use FILL  FILL_5001
timestamp 1018054153
transform 1 0 7200 0 1 4480
box -16 -6 32 210
use FILL  FILL_5003
timestamp 1018054153
transform 1 0 7216 0 1 4480
box -16 -6 32 210
use FILL  FILL_5005
timestamp 1018054153
transform 1 0 7232 0 1 4480
box -16 -6 32 210
use FILL  FILL_5007
timestamp 1018054153
transform 1 0 7248 0 1 4480
box -16 -6 32 210
use FILL  FILL_5009
timestamp 1018054153
transform 1 0 7264 0 1 4480
box -16 -6 32 210
use FILL  FILL_5011
timestamp 1018054153
transform 1 0 7280 0 1 4480
box -16 -6 32 210
use FILL  FILL_5013
timestamp 1018054153
transform 1 0 7296 0 1 4480
box -16 -6 32 210
use FILL  FILL_5015
timestamp 1018054153
transform 1 0 7312 0 1 4480
box -16 -6 32 210
use FILL  FILL_5017
timestamp 1018054153
transform 1 0 7328 0 1 4480
box -16 -6 32 210
use FILL  FILL_5019
timestamp 1018054153
transform 1 0 7344 0 1 4480
box -16 -6 32 210
use FILL  FILL_5021
timestamp 1018054153
transform 1 0 7360 0 1 4480
box -16 -6 32 210
use FILL  FILL_5023
timestamp 1018054153
transform 1 0 7376 0 1 4480
box -16 -6 32 210
use FILL  FILL_5025
timestamp 1018054153
transform 1 0 7392 0 1 4480
box -16 -6 32 210
use FILL  FILL_5027
timestamp 1018054153
transform 1 0 7408 0 1 4480
box -16 -6 32 210
use FILL  FILL_5029
timestamp 1018054153
transform 1 0 7424 0 1 4480
box -16 -6 32 210
use FILL  FILL_5031
timestamp 1018054153
transform 1 0 7440 0 1 4480
box -16 -6 32 210
use FILL  FILL_5033
timestamp 1018054153
transform 1 0 7456 0 1 4480
box -16 -6 32 210
use FILL  FILL_5035
timestamp 1018054153
transform 1 0 7472 0 1 4480
box -16 -6 32 210
use FILL  FILL_5037
timestamp 1018054153
transform 1 0 7488 0 1 4480
box -16 -6 32 210
use FILL  FILL_5039
timestamp 1018054153
transform 1 0 7504 0 1 4480
box -16 -6 32 210
use FILL  FILL_5041
timestamp 1018054153
transform 1 0 7520 0 1 4480
box -16 -6 32 210
use FILL  FILL_5043
timestamp 1018054153
transform 1 0 7536 0 1 4480
box -16 -6 32 210
use FILL  FILL_5045
timestamp 1018054153
transform 1 0 7552 0 1 4480
box -16 -6 32 210
use FILL  FILL_5047
timestamp 1018054153
transform 1 0 7568 0 1 4480
box -16 -6 32 210
use FILL  FILL_5049
timestamp 1018054153
transform 1 0 7584 0 1 4480
box -16 -6 32 210
use FILL  FILL_5051
timestamp 1018054153
transform 1 0 7600 0 1 4480
box -16 -6 32 210
use FILL  FILL_5053
timestamp 1018054153
transform 1 0 7616 0 1 4480
box -16 -6 32 210
use FILL  FILL_5055
timestamp 1018054153
transform 1 0 7632 0 1 4480
box -16 -6 32 210
use FILL  FILL_5057
timestamp 1018054153
transform 1 0 7648 0 1 4480
box -16 -6 32 210
use FILL  FILL_5059
timestamp 1018054153
transform 1 0 7664 0 1 4480
box -16 -6 32 210
use FILL  FILL_5061
timestamp 1018054153
transform 1 0 7680 0 1 4480
box -16 -6 32 210
use FILL  FILL_5063
timestamp 1018054153
transform 1 0 7696 0 1 4480
box -16 -6 32 210
use FILL  FILL_5065
timestamp 1018054153
transform 1 0 7712 0 1 4480
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_29
timestamp 1542725905
transform 1 0 7908 0 1 4480
box -48 -6 48 6
use M2_M1  M2_M1_242
timestamp 1542725905
transform 1 0 6872 0 1 4410
box -4 -4 4 4
use M2_M1  M2_M1_243
timestamp 1542725905
transform 1 0 7672 0 1 4410
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_30
timestamp 1542725905
transform 1 0 2212 0 1 4280
box -48 -6 48 6
use FILL  FILL_4601
timestamp 1018054153
transform 1 0 2272 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4603
timestamp 1018054153
transform 1 0 2288 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4605
timestamp 1018054153
transform 1 0 2304 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4607
timestamp 1018054153
transform 1 0 2320 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4609
timestamp 1018054153
transform 1 0 2336 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4611
timestamp 1018054153
transform 1 0 2352 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4613
timestamp 1018054153
transform 1 0 2368 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4615
timestamp 1018054153
transform 1 0 2384 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4617
timestamp 1018054153
transform 1 0 2400 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4619
timestamp 1018054153
transform 1 0 2416 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4621
timestamp 1018054153
transform 1 0 2432 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4623
timestamp 1018054153
transform 1 0 2448 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4625
timestamp 1018054153
transform 1 0 2464 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4627
timestamp 1018054153
transform 1 0 2480 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4629
timestamp 1018054153
transform 1 0 2496 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4631
timestamp 1018054153
transform 1 0 2512 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4633
timestamp 1018054153
transform 1 0 2528 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4635
timestamp 1018054153
transform 1 0 2544 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4637
timestamp 1018054153
transform 1 0 2560 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4639
timestamp 1018054153
transform 1 0 2576 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4641
timestamp 1018054153
transform 1 0 2592 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4643
timestamp 1018054153
transform 1 0 2608 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4645
timestamp 1018054153
transform 1 0 2624 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4647
timestamp 1018054153
transform 1 0 2640 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4649
timestamp 1018054153
transform 1 0 2656 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4651
timestamp 1018054153
transform 1 0 2672 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4653
timestamp 1018054153
transform 1 0 2688 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4655
timestamp 1018054153
transform 1 0 2704 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4657
timestamp 1018054153
transform 1 0 2720 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4659
timestamp 1018054153
transform 1 0 2736 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4661
timestamp 1018054153
transform 1 0 2752 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4663
timestamp 1018054153
transform 1 0 2768 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4665
timestamp 1018054153
transform 1 0 2784 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4667
timestamp 1018054153
transform 1 0 2800 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4669
timestamp 1018054153
transform 1 0 2816 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4671
timestamp 1018054153
transform 1 0 2832 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4673
timestamp 1018054153
transform 1 0 2848 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4675
timestamp 1018054153
transform 1 0 2864 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4677
timestamp 1018054153
transform 1 0 2880 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4679
timestamp 1018054153
transform 1 0 2896 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4681
timestamp 1018054153
transform 1 0 2912 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4683
timestamp 1018054153
transform 1 0 2928 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4685
timestamp 1018054153
transform 1 0 2944 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4687
timestamp 1018054153
transform 1 0 2960 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4689
timestamp 1018054153
transform 1 0 2976 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4691
timestamp 1018054153
transform 1 0 2992 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4693
timestamp 1018054153
transform 1 0 3008 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4695
timestamp 1018054153
transform 1 0 3024 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4697
timestamp 1018054153
transform 1 0 3040 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4699
timestamp 1018054153
transform 1 0 3056 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4701
timestamp 1018054153
transform 1 0 3072 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4703
timestamp 1018054153
transform 1 0 3088 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4705
timestamp 1018054153
transform 1 0 3104 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4707
timestamp 1018054153
transform 1 0 3120 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4709
timestamp 1018054153
transform 1 0 3136 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4711
timestamp 1018054153
transform 1 0 3152 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4713
timestamp 1018054153
transform 1 0 3168 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4715
timestamp 1018054153
transform 1 0 3184 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4717
timestamp 1018054153
transform 1 0 3200 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4719
timestamp 1018054153
transform 1 0 3216 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4721
timestamp 1018054153
transform 1 0 3232 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4723
timestamp 1018054153
transform 1 0 3248 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4725
timestamp 1018054153
transform 1 0 3264 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4727
timestamp 1018054153
transform 1 0 3280 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4729
timestamp 1018054153
transform 1 0 3296 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4731
timestamp 1018054153
transform 1 0 3312 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4733
timestamp 1018054153
transform 1 0 3328 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4735
timestamp 1018054153
transform 1 0 3344 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4737
timestamp 1018054153
transform 1 0 3360 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4739
timestamp 1018054153
transform 1 0 3376 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4741
timestamp 1018054153
transform 1 0 3392 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4743
timestamp 1018054153
transform 1 0 3408 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4745
timestamp 1018054153
transform 1 0 3424 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4747
timestamp 1018054153
transform 1 0 3440 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4749
timestamp 1018054153
transform 1 0 3456 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4751
timestamp 1018054153
transform 1 0 3472 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4753
timestamp 1018054153
transform 1 0 3488 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4755
timestamp 1018054153
transform 1 0 3504 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4757
timestamp 1018054153
transform 1 0 3520 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4759
timestamp 1018054153
transform 1 0 3536 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4761
timestamp 1018054153
transform 1 0 3552 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4763
timestamp 1018054153
transform 1 0 3568 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4765
timestamp 1018054153
transform 1 0 3584 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4767
timestamp 1018054153
transform 1 0 3600 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4769
timestamp 1018054153
transform 1 0 3616 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4771
timestamp 1018054153
transform 1 0 3632 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4773
timestamp 1018054153
transform 1 0 3648 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4775
timestamp 1018054153
transform 1 0 3664 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4777
timestamp 1018054153
transform 1 0 3680 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4779
timestamp 1018054153
transform 1 0 3696 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4781
timestamp 1018054153
transform 1 0 3712 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4783
timestamp 1018054153
transform 1 0 3728 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4785
timestamp 1018054153
transform 1 0 3744 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4787
timestamp 1018054153
transform 1 0 3760 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4789
timestamp 1018054153
transform 1 0 3776 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4790
timestamp 1018054153
transform 1 0 3792 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4791
timestamp 1018054153
transform 1 0 3808 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4792
timestamp 1018054153
transform 1 0 3824 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4793
timestamp 1018054153
transform 1 0 3840 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4794
timestamp 1018054153
transform 1 0 3856 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4795
timestamp 1018054153
transform 1 0 3872 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4796
timestamp 1018054153
transform 1 0 3888 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4797
timestamp 1018054153
transform 1 0 3904 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4798
timestamp 1018054153
transform 1 0 3920 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4799
timestamp 1018054153
transform 1 0 3936 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4800
timestamp 1018054153
transform 1 0 3952 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4801
timestamp 1018054153
transform 1 0 3968 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4802
timestamp 1018054153
transform 1 0 3984 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4803
timestamp 1018054153
transform 1 0 4000 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4804
timestamp 1018054153
transform 1 0 4016 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4805
timestamp 1018054153
transform 1 0 4032 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4806
timestamp 1018054153
transform 1 0 4048 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4807
timestamp 1018054153
transform 1 0 4064 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4808
timestamp 1018054153
transform 1 0 4080 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4809
timestamp 1018054153
transform 1 0 4096 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4810
timestamp 1018054153
transform 1 0 4112 0 -1 4480
box -16 -6 32 210
use M3_M2  M3_M2_98
timestamp 1542725905
transform 1 0 4152 0 1 4290
box -6 -6 6 6
use FILL  FILL_4811
timestamp 1018054153
transform 1 0 4128 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4813
timestamp 1018054153
transform 1 0 4144 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4815
timestamp 1018054153
transform 1 0 4160 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4817
timestamp 1018054153
transform 1 0 4176 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4819
timestamp 1018054153
transform 1 0 4192 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4821
timestamp 1018054153
transform 1 0 4208 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4823
timestamp 1018054153
transform 1 0 4224 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4825
timestamp 1018054153
transform 1 0 4240 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4827
timestamp 1018054153
transform 1 0 4256 0 -1 4480
box -16 -6 32 210
use M2_M1  M2_M1_252
timestamp 1542725905
transform 1 0 4296 0 1 4280
box -4 -4 4 4
use M3_M2  M3_M2_99
timestamp 1542725905
transform 1 0 4440 0 1 4290
box -6 -6 6 6
use DFFSR  DFFSR_1
timestamp 1071163401
transform 1 0 4272 0 -1 4480
box -16 -6 368 210
use FILL  FILL_4850
timestamp 1018054153
transform 1 0 4624 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4851
timestamp 1018054153
transform 1 0 4640 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4852
timestamp 1018054153
transform 1 0 4656 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4853
timestamp 1018054153
transform 1 0 4672 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4854
timestamp 1018054153
transform 1 0 4688 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4855
timestamp 1018054153
transform 1 0 4704 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4856
timestamp 1018054153
transform 1 0 4720 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4857
timestamp 1018054153
transform 1 0 4736 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4858
timestamp 1018054153
transform 1 0 4752 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4859
timestamp 1018054153
transform 1 0 4768 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4860
timestamp 1018054153
transform 1 0 4784 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4861
timestamp 1018054153
transform 1 0 4800 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4862
timestamp 1018054153
transform 1 0 4816 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4863
timestamp 1018054153
transform 1 0 4832 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4864
timestamp 1018054153
transform 1 0 4848 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4865
timestamp 1018054153
transform 1 0 4864 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4866
timestamp 1018054153
transform 1 0 4880 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4867
timestamp 1018054153
transform 1 0 4896 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4868
timestamp 1018054153
transform 1 0 4912 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4869
timestamp 1018054153
transform 1 0 4928 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4870
timestamp 1018054153
transform 1 0 4944 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4871
timestamp 1018054153
transform 1 0 4960 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4872
timestamp 1018054153
transform 1 0 4976 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4873
timestamp 1018054153
transform 1 0 4992 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4874
timestamp 1018054153
transform 1 0 5008 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4875
timestamp 1018054153
transform 1 0 5024 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4876
timestamp 1018054153
transform 1 0 5040 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4877
timestamp 1018054153
transform 1 0 5056 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4878
timestamp 1018054153
transform 1 0 5072 0 -1 4480
box -16 -6 32 210
use M2_M1  M2_M1_253
timestamp 1542725905
transform 1 0 5128 0 1 4280
box -4 -4 4 4
use M3_M2  M3_M2_100
timestamp 1542725905
transform 1 0 5176 0 1 4290
box -6 -6 6 6
use M3_M2  M3_M2_101
timestamp 1542725905
transform 1 0 5256 0 1 4290
box -6 -6 6 6
use M2_M1  M2_M1_254
timestamp 1542725905
transform 1 0 5416 0 1 4280
box -4 -4 4 4
use DFFSR  DFFSR_2
timestamp 1071163401
transform 1 0 5088 0 -1 4480
box -16 -6 368 210
use FILL  FILL_4879
timestamp 1018054153
transform 1 0 5440 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4880
timestamp 1018054153
transform 1 0 5456 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4881
timestamp 1018054153
transform 1 0 5472 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4882
timestamp 1018054153
transform 1 0 5488 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4883
timestamp 1018054153
transform 1 0 5504 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4884
timestamp 1018054153
transform 1 0 5520 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4885
timestamp 1018054153
transform 1 0 5536 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4886
timestamp 1018054153
transform 1 0 5552 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4887
timestamp 1018054153
transform 1 0 5568 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4888
timestamp 1018054153
transform 1 0 5584 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4889
timestamp 1018054153
transform 1 0 5600 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4890
timestamp 1018054153
transform 1 0 5616 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4891
timestamp 1018054153
transform 1 0 5632 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4892
timestamp 1018054153
transform 1 0 5648 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4893
timestamp 1018054153
transform 1 0 5664 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4894
timestamp 1018054153
transform 1 0 5680 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4895
timestamp 1018054153
transform 1 0 5696 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4896
timestamp 1018054153
transform 1 0 5712 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4897
timestamp 1018054153
transform 1 0 5728 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4898
timestamp 1018054153
transform 1 0 5744 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4899
timestamp 1018054153
transform 1 0 5760 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4900
timestamp 1018054153
transform 1 0 5776 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4901
timestamp 1018054153
transform 1 0 5792 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4902
timestamp 1018054153
transform 1 0 5808 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4903
timestamp 1018054153
transform 1 0 5824 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4904
timestamp 1018054153
transform 1 0 5840 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4905
timestamp 1018054153
transform 1 0 5856 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4906
timestamp 1018054153
transform 1 0 5872 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4907
timestamp 1018054153
transform 1 0 5888 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4908
timestamp 1018054153
transform 1 0 5904 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4909
timestamp 1018054153
transform 1 0 5920 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4910
timestamp 1018054153
transform 1 0 5936 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4911
timestamp 1018054153
transform 1 0 5952 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4912
timestamp 1018054153
transform 1 0 5968 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4913
timestamp 1018054153
transform 1 0 5984 0 -1 4480
box -16 -6 32 210
use M2_M1  M2_M1_255
timestamp 1542725905
transform 1 0 6040 0 1 4280
box -4 -4 4 4
use DFFSR  DFFSR_3
timestamp 1071163401
transform 1 0 6000 0 -1 4480
box -16 -6 368 210
use FILL  FILL_4914
timestamp 1018054153
transform 1 0 6352 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4915
timestamp 1018054153
transform 1 0 6368 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4916
timestamp 1018054153
transform 1 0 6384 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4917
timestamp 1018054153
transform 1 0 6400 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4918
timestamp 1018054153
transform 1 0 6416 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4919
timestamp 1018054153
transform 1 0 6432 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4920
timestamp 1018054153
transform 1 0 6448 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4921
timestamp 1018054153
transform 1 0 6464 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4922
timestamp 1018054153
transform 1 0 6480 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4923
timestamp 1018054153
transform 1 0 6496 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4924
timestamp 1018054153
transform 1 0 6512 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4925
timestamp 1018054153
transform 1 0 6528 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4926
timestamp 1018054153
transform 1 0 6544 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4927
timestamp 1018054153
transform 1 0 6560 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4928
timestamp 1018054153
transform 1 0 6576 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4929
timestamp 1018054153
transform 1 0 6592 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4931
timestamp 1018054153
transform 1 0 6608 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4933
timestamp 1018054153
transform 1 0 6624 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4935
timestamp 1018054153
transform 1 0 6640 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4937
timestamp 1018054153
transform 1 0 6656 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4939
timestamp 1018054153
transform 1 0 6672 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4941
timestamp 1018054153
transform 1 0 6688 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4943
timestamp 1018054153
transform 1 0 6704 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4945
timestamp 1018054153
transform 1 0 6720 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4947
timestamp 1018054153
transform 1 0 6736 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4949
timestamp 1018054153
transform 1 0 6752 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4951
timestamp 1018054153
transform 1 0 6768 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4953
timestamp 1018054153
transform 1 0 6784 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4955
timestamp 1018054153
transform 1 0 6800 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4957
timestamp 1018054153
transform 1 0 6816 0 -1 4480
box -16 -6 32 210
use BUFX2  BUFX2_2
timestamp 1090542073
transform 1 0 6832 0 -1 4480
box -10 -6 56 210
use FILL  FILL_4962
timestamp 1018054153
transform 1 0 6880 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4964
timestamp 1018054153
transform 1 0 6896 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4966
timestamp 1018054153
transform 1 0 6912 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4968
timestamp 1018054153
transform 1 0 6928 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4970
timestamp 1018054153
transform 1 0 6944 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4972
timestamp 1018054153
transform 1 0 6960 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4974
timestamp 1018054153
transform 1 0 6976 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4976
timestamp 1018054153
transform 1 0 6992 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4978
timestamp 1018054153
transform 1 0 7008 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4980
timestamp 1018054153
transform 1 0 7024 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4982
timestamp 1018054153
transform 1 0 7040 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4984
timestamp 1018054153
transform 1 0 7056 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4986
timestamp 1018054153
transform 1 0 7072 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4988
timestamp 1018054153
transform 1 0 7088 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4990
timestamp 1018054153
transform 1 0 7104 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4992
timestamp 1018054153
transform 1 0 7120 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4994
timestamp 1018054153
transform 1 0 7136 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4996
timestamp 1018054153
transform 1 0 7152 0 -1 4480
box -16 -6 32 210
use FILL  FILL_4998
timestamp 1018054153
transform 1 0 7168 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5000
timestamp 1018054153
transform 1 0 7184 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5002
timestamp 1018054153
transform 1 0 7200 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5004
timestamp 1018054153
transform 1 0 7216 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5006
timestamp 1018054153
transform 1 0 7232 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5008
timestamp 1018054153
transform 1 0 7248 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5010
timestamp 1018054153
transform 1 0 7264 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5012
timestamp 1018054153
transform 1 0 7280 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5014
timestamp 1018054153
transform 1 0 7296 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5016
timestamp 1018054153
transform 1 0 7312 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5018
timestamp 1018054153
transform 1 0 7328 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5020
timestamp 1018054153
transform 1 0 7344 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5022
timestamp 1018054153
transform 1 0 7360 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5024
timestamp 1018054153
transform 1 0 7376 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5026
timestamp 1018054153
transform 1 0 7392 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5028
timestamp 1018054153
transform 1 0 7408 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5030
timestamp 1018054153
transform 1 0 7424 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5032
timestamp 1018054153
transform 1 0 7440 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5034
timestamp 1018054153
transform 1 0 7456 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5036
timestamp 1018054153
transform 1 0 7472 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5038
timestamp 1018054153
transform 1 0 7488 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5040
timestamp 1018054153
transform 1 0 7504 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5042
timestamp 1018054153
transform 1 0 7520 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5044
timestamp 1018054153
transform 1 0 7536 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5046
timestamp 1018054153
transform 1 0 7552 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5048
timestamp 1018054153
transform 1 0 7568 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5050
timestamp 1018054153
transform 1 0 7584 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5052
timestamp 1018054153
transform 1 0 7600 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5054
timestamp 1018054153
transform 1 0 7616 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5056
timestamp 1018054153
transform 1 0 7632 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5058
timestamp 1018054153
transform 1 0 7648 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5060
timestamp 1018054153
transform 1 0 7664 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5062
timestamp 1018054153
transform 1 0 7680 0 -1 4480
box -16 -6 32 210
use FILL  FILL_5064
timestamp 1018054153
transform 1 0 7696 0 -1 4480
box -16 -6 32 210
use PADOUT  PADOUT_1
timestamp 1084294529
transform 0 1 8000 -1 0 5000
box -12 -6 606 2000
use M3_M2  M3_M2_97
timestamp 1542725905
transform 1 0 8002 0 1 4310
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_31
timestamp 1542725905
transform 1 0 7788 0 1 4280
box -48 -6 48 6
use FILL  FILL_5066
timestamp 1018054153
transform 1 0 7712 0 -1 4480
box -16 -6 32 210
use M3_M2  M3_M2_102
timestamp 1542725905
transform 1 0 5112 0 1 4190
box -6 -6 6 6
use M3_M2  M3_M2_105
timestamp 1542725905
transform 1 0 5176 0 1 4130
box -6 -6 6 6
use M3_M2  M3_M2_106
timestamp 1542725905
transform 1 0 5208 0 1 4130
box -6 -6 6 6
use M2_M1  M2_M1_256
timestamp 1542725905
transform 1 0 5416 0 1 4190
box -4 -4 4 4
use M3_M2  M3_M2_103
timestamp 1542725905
transform 1 0 5464 0 1 4190
box -6 -6 6 6
use M2_M1  M2_M1_257
timestamp 1542725905
transform 1 0 5464 0 1 4170
box -4 -4 4 4
use M2_M1  M2_M1_258
timestamp 1542725905
transform 1 0 5528 0 1 4150
box -4 -4 4 4
use M3_M2  M3_M2_107
timestamp 1542725905
transform 1 0 5528 0 1 4130
box -6 -6 6 6
use M2_M1  M2_M1_260
timestamp 1542725905
transform 1 0 5560 0 1 4126
box -4 -4 4 4
use M3_M2  M3_M2_104
timestamp 1542725905
transform 1 0 5880 0 1 4190
box -6 -6 6 6
use M3_M2  M3_M2_108
timestamp 1542725905
transform 1 0 5976 0 1 4130
box -6 -6 6 6
use M3_M2  M3_M2_109
timestamp 1542725905
transform 1 0 6168 0 1 4130
box -6 -6 6 6
use M2_M1  M2_M1_259
timestamp 1542725905
transform 1 0 6280 0 1 4150
box -4 -4 4 4
use M3_M2  M3_M2_110
timestamp 1542725905
transform 1 0 6952 0 1 4130
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_32
timestamp 1542725905
transform 1 0 2092 0 1 4080
box -48 -6 48 6
use FILL  FILL_5067
timestamp 1018054153
transform 1 0 2272 0 1 4080
box -16 -6 32 210
use FILL  FILL_5069
timestamp 1018054153
transform 1 0 2288 0 1 4080
box -16 -6 32 210
use FILL  FILL_5071
timestamp 1018054153
transform 1 0 2304 0 1 4080
box -16 -6 32 210
use FILL  FILL_5073
timestamp 1018054153
transform 1 0 2320 0 1 4080
box -16 -6 32 210
use FILL  FILL_5075
timestamp 1018054153
transform 1 0 2336 0 1 4080
box -16 -6 32 210
use FILL  FILL_5077
timestamp 1018054153
transform 1 0 2352 0 1 4080
box -16 -6 32 210
use FILL  FILL_5079
timestamp 1018054153
transform 1 0 2368 0 1 4080
box -16 -6 32 210
use FILL  FILL_5081
timestamp 1018054153
transform 1 0 2384 0 1 4080
box -16 -6 32 210
use FILL  FILL_5083
timestamp 1018054153
transform 1 0 2400 0 1 4080
box -16 -6 32 210
use FILL  FILL_5085
timestamp 1018054153
transform 1 0 2416 0 1 4080
box -16 -6 32 210
use FILL  FILL_5087
timestamp 1018054153
transform 1 0 2432 0 1 4080
box -16 -6 32 210
use FILL  FILL_5089
timestamp 1018054153
transform 1 0 2448 0 1 4080
box -16 -6 32 210
use FILL  FILL_5091
timestamp 1018054153
transform 1 0 2464 0 1 4080
box -16 -6 32 210
use FILL  FILL_5093
timestamp 1018054153
transform 1 0 2480 0 1 4080
box -16 -6 32 210
use FILL  FILL_5095
timestamp 1018054153
transform 1 0 2496 0 1 4080
box -16 -6 32 210
use FILL  FILL_5097
timestamp 1018054153
transform 1 0 2512 0 1 4080
box -16 -6 32 210
use FILL  FILL_5099
timestamp 1018054153
transform 1 0 2528 0 1 4080
box -16 -6 32 210
use FILL  FILL_5101
timestamp 1018054153
transform 1 0 2544 0 1 4080
box -16 -6 32 210
use FILL  FILL_5103
timestamp 1018054153
transform 1 0 2560 0 1 4080
box -16 -6 32 210
use FILL  FILL_5105
timestamp 1018054153
transform 1 0 2576 0 1 4080
box -16 -6 32 210
use FILL  FILL_5107
timestamp 1018054153
transform 1 0 2592 0 1 4080
box -16 -6 32 210
use FILL  FILL_5109
timestamp 1018054153
transform 1 0 2608 0 1 4080
box -16 -6 32 210
use FILL  FILL_5111
timestamp 1018054153
transform 1 0 2624 0 1 4080
box -16 -6 32 210
use FILL  FILL_5113
timestamp 1018054153
transform 1 0 2640 0 1 4080
box -16 -6 32 210
use FILL  FILL_5115
timestamp 1018054153
transform 1 0 2656 0 1 4080
box -16 -6 32 210
use FILL  FILL_5117
timestamp 1018054153
transform 1 0 2672 0 1 4080
box -16 -6 32 210
use FILL  FILL_5119
timestamp 1018054153
transform 1 0 2688 0 1 4080
box -16 -6 32 210
use FILL  FILL_5121
timestamp 1018054153
transform 1 0 2704 0 1 4080
box -16 -6 32 210
use FILL  FILL_5123
timestamp 1018054153
transform 1 0 2720 0 1 4080
box -16 -6 32 210
use FILL  FILL_5125
timestamp 1018054153
transform 1 0 2736 0 1 4080
box -16 -6 32 210
use FILL  FILL_5127
timestamp 1018054153
transform 1 0 2752 0 1 4080
box -16 -6 32 210
use FILL  FILL_5129
timestamp 1018054153
transform 1 0 2768 0 1 4080
box -16 -6 32 210
use FILL  FILL_5131
timestamp 1018054153
transform 1 0 2784 0 1 4080
box -16 -6 32 210
use FILL  FILL_5133
timestamp 1018054153
transform 1 0 2800 0 1 4080
box -16 -6 32 210
use FILL  FILL_5135
timestamp 1018054153
transform 1 0 2816 0 1 4080
box -16 -6 32 210
use FILL  FILL_5137
timestamp 1018054153
transform 1 0 2832 0 1 4080
box -16 -6 32 210
use FILL  FILL_5139
timestamp 1018054153
transform 1 0 2848 0 1 4080
box -16 -6 32 210
use FILL  FILL_5141
timestamp 1018054153
transform 1 0 2864 0 1 4080
box -16 -6 32 210
use FILL  FILL_5143
timestamp 1018054153
transform 1 0 2880 0 1 4080
box -16 -6 32 210
use FILL  FILL_5145
timestamp 1018054153
transform 1 0 2896 0 1 4080
box -16 -6 32 210
use FILL  FILL_5147
timestamp 1018054153
transform 1 0 2912 0 1 4080
box -16 -6 32 210
use FILL  FILL_5149
timestamp 1018054153
transform 1 0 2928 0 1 4080
box -16 -6 32 210
use FILL  FILL_5151
timestamp 1018054153
transform 1 0 2944 0 1 4080
box -16 -6 32 210
use FILL  FILL_5153
timestamp 1018054153
transform 1 0 2960 0 1 4080
box -16 -6 32 210
use FILL  FILL_5155
timestamp 1018054153
transform 1 0 2976 0 1 4080
box -16 -6 32 210
use FILL  FILL_5157
timestamp 1018054153
transform 1 0 2992 0 1 4080
box -16 -6 32 210
use FILL  FILL_5159
timestamp 1018054153
transform 1 0 3008 0 1 4080
box -16 -6 32 210
use FILL  FILL_5161
timestamp 1018054153
transform 1 0 3024 0 1 4080
box -16 -6 32 210
use FILL  FILL_5163
timestamp 1018054153
transform 1 0 3040 0 1 4080
box -16 -6 32 210
use FILL  FILL_5165
timestamp 1018054153
transform 1 0 3056 0 1 4080
box -16 -6 32 210
use FILL  FILL_5167
timestamp 1018054153
transform 1 0 3072 0 1 4080
box -16 -6 32 210
use FILL  FILL_5169
timestamp 1018054153
transform 1 0 3088 0 1 4080
box -16 -6 32 210
use FILL  FILL_5171
timestamp 1018054153
transform 1 0 3104 0 1 4080
box -16 -6 32 210
use FILL  FILL_5173
timestamp 1018054153
transform 1 0 3120 0 1 4080
box -16 -6 32 210
use FILL  FILL_5175
timestamp 1018054153
transform 1 0 3136 0 1 4080
box -16 -6 32 210
use FILL  FILL_5177
timestamp 1018054153
transform 1 0 3152 0 1 4080
box -16 -6 32 210
use FILL  FILL_5179
timestamp 1018054153
transform 1 0 3168 0 1 4080
box -16 -6 32 210
use FILL  FILL_5181
timestamp 1018054153
transform 1 0 3184 0 1 4080
box -16 -6 32 210
use FILL  FILL_5183
timestamp 1018054153
transform 1 0 3200 0 1 4080
box -16 -6 32 210
use FILL  FILL_5185
timestamp 1018054153
transform 1 0 3216 0 1 4080
box -16 -6 32 210
use FILL  FILL_5187
timestamp 1018054153
transform 1 0 3232 0 1 4080
box -16 -6 32 210
use FILL  FILL_5189
timestamp 1018054153
transform 1 0 3248 0 1 4080
box -16 -6 32 210
use FILL  FILL_5191
timestamp 1018054153
transform 1 0 3264 0 1 4080
box -16 -6 32 210
use FILL  FILL_5193
timestamp 1018054153
transform 1 0 3280 0 1 4080
box -16 -6 32 210
use FILL  FILL_5195
timestamp 1018054153
transform 1 0 3296 0 1 4080
box -16 -6 32 210
use FILL  FILL_5197
timestamp 1018054153
transform 1 0 3312 0 1 4080
box -16 -6 32 210
use FILL  FILL_5199
timestamp 1018054153
transform 1 0 3328 0 1 4080
box -16 -6 32 210
use FILL  FILL_5201
timestamp 1018054153
transform 1 0 3344 0 1 4080
box -16 -6 32 210
use FILL  FILL_5203
timestamp 1018054153
transform 1 0 3360 0 1 4080
box -16 -6 32 210
use FILL  FILL_5205
timestamp 1018054153
transform 1 0 3376 0 1 4080
box -16 -6 32 210
use FILL  FILL_5207
timestamp 1018054153
transform 1 0 3392 0 1 4080
box -16 -6 32 210
use FILL  FILL_5209
timestamp 1018054153
transform 1 0 3408 0 1 4080
box -16 -6 32 210
use FILL  FILL_5211
timestamp 1018054153
transform 1 0 3424 0 1 4080
box -16 -6 32 210
use FILL  FILL_5213
timestamp 1018054153
transform 1 0 3440 0 1 4080
box -16 -6 32 210
use FILL  FILL_5215
timestamp 1018054153
transform 1 0 3456 0 1 4080
box -16 -6 32 210
use FILL  FILL_5217
timestamp 1018054153
transform 1 0 3472 0 1 4080
box -16 -6 32 210
use FILL  FILL_5219
timestamp 1018054153
transform 1 0 3488 0 1 4080
box -16 -6 32 210
use FILL  FILL_5221
timestamp 1018054153
transform 1 0 3504 0 1 4080
box -16 -6 32 210
use FILL  FILL_5223
timestamp 1018054153
transform 1 0 3520 0 1 4080
box -16 -6 32 210
use FILL  FILL_5225
timestamp 1018054153
transform 1 0 3536 0 1 4080
box -16 -6 32 210
use FILL  FILL_5227
timestamp 1018054153
transform 1 0 3552 0 1 4080
box -16 -6 32 210
use FILL  FILL_5229
timestamp 1018054153
transform 1 0 3568 0 1 4080
box -16 -6 32 210
use FILL  FILL_5231
timestamp 1018054153
transform 1 0 3584 0 1 4080
box -16 -6 32 210
use FILL  FILL_5233
timestamp 1018054153
transform 1 0 3600 0 1 4080
box -16 -6 32 210
use FILL  FILL_5235
timestamp 1018054153
transform 1 0 3616 0 1 4080
box -16 -6 32 210
use FILL  FILL_5237
timestamp 1018054153
transform 1 0 3632 0 1 4080
box -16 -6 32 210
use FILL  FILL_5239
timestamp 1018054153
transform 1 0 3648 0 1 4080
box -16 -6 32 210
use FILL  FILL_5241
timestamp 1018054153
transform 1 0 3664 0 1 4080
box -16 -6 32 210
use FILL  FILL_5243
timestamp 1018054153
transform 1 0 3680 0 1 4080
box -16 -6 32 210
use FILL  FILL_5245
timestamp 1018054153
transform 1 0 3696 0 1 4080
box -16 -6 32 210
use FILL  FILL_5247
timestamp 1018054153
transform 1 0 3712 0 1 4080
box -16 -6 32 210
use FILL  FILL_5249
timestamp 1018054153
transform 1 0 3728 0 1 4080
box -16 -6 32 210
use FILL  FILL_5251
timestamp 1018054153
transform 1 0 3744 0 1 4080
box -16 -6 32 210
use FILL  FILL_5253
timestamp 1018054153
transform 1 0 3760 0 1 4080
box -16 -6 32 210
use FILL  FILL_5255
timestamp 1018054153
transform 1 0 3776 0 1 4080
box -16 -6 32 210
use FILL  FILL_5257
timestamp 1018054153
transform 1 0 3792 0 1 4080
box -16 -6 32 210
use FILL  FILL_5259
timestamp 1018054153
transform 1 0 3808 0 1 4080
box -16 -6 32 210
use FILL  FILL_5261
timestamp 1018054153
transform 1 0 3824 0 1 4080
box -16 -6 32 210
use FILL  FILL_5263
timestamp 1018054153
transform 1 0 3840 0 1 4080
box -16 -6 32 210
use FILL  FILL_5265
timestamp 1018054153
transform 1 0 3856 0 1 4080
box -16 -6 32 210
use FILL  FILL_5267
timestamp 1018054153
transform 1 0 3872 0 1 4080
box -16 -6 32 210
use FILL  FILL_5269
timestamp 1018054153
transform 1 0 3888 0 1 4080
box -16 -6 32 210
use FILL  FILL_5271
timestamp 1018054153
transform 1 0 3904 0 1 4080
box -16 -6 32 210
use FILL  FILL_5273
timestamp 1018054153
transform 1 0 3920 0 1 4080
box -16 -6 32 210
use FILL  FILL_5275
timestamp 1018054153
transform 1 0 3936 0 1 4080
box -16 -6 32 210
use FILL  FILL_5277
timestamp 1018054153
transform 1 0 3952 0 1 4080
box -16 -6 32 210
use FILL  FILL_5279
timestamp 1018054153
transform 1 0 3968 0 1 4080
box -16 -6 32 210
use FILL  FILL_5281
timestamp 1018054153
transform 1 0 3984 0 1 4080
box -16 -6 32 210
use FILL  FILL_5283
timestamp 1018054153
transform 1 0 4000 0 1 4080
box -16 -6 32 210
use FILL  FILL_5285
timestamp 1018054153
transform 1 0 4016 0 1 4080
box -16 -6 32 210
use FILL  FILL_5287
timestamp 1018054153
transform 1 0 4032 0 1 4080
box -16 -6 32 210
use FILL  FILL_5289
timestamp 1018054153
transform 1 0 4048 0 1 4080
box -16 -6 32 210
use FILL  FILL_5291
timestamp 1018054153
transform 1 0 4064 0 1 4080
box -16 -6 32 210
use FILL  FILL_5293
timestamp 1018054153
transform 1 0 4080 0 1 4080
box -16 -6 32 210
use FILL  FILL_5295
timestamp 1018054153
transform 1 0 4096 0 1 4080
box -16 -6 32 210
use FILL  FILL_5297
timestamp 1018054153
transform 1 0 4112 0 1 4080
box -16 -6 32 210
use FILL  FILL_5299
timestamp 1018054153
transform 1 0 4128 0 1 4080
box -16 -6 32 210
use FILL  FILL_5301
timestamp 1018054153
transform 1 0 4144 0 1 4080
box -16 -6 32 210
use FILL  FILL_5303
timestamp 1018054153
transform 1 0 4160 0 1 4080
box -16 -6 32 210
use FILL  FILL_5305
timestamp 1018054153
transform 1 0 4176 0 1 4080
box -16 -6 32 210
use FILL  FILL_5307
timestamp 1018054153
transform 1 0 4192 0 1 4080
box -16 -6 32 210
use FILL  FILL_5309
timestamp 1018054153
transform 1 0 4208 0 1 4080
box -16 -6 32 210
use FILL  FILL_5311
timestamp 1018054153
transform 1 0 4224 0 1 4080
box -16 -6 32 210
use FILL  FILL_5313
timestamp 1018054153
transform 1 0 4240 0 1 4080
box -16 -6 32 210
use FILL  FILL_5315
timestamp 1018054153
transform 1 0 4256 0 1 4080
box -16 -6 32 210
use FILL  FILL_5317
timestamp 1018054153
transform 1 0 4272 0 1 4080
box -16 -6 32 210
use FILL  FILL_5319
timestamp 1018054153
transform 1 0 4288 0 1 4080
box -16 -6 32 210
use FILL  FILL_5321
timestamp 1018054153
transform 1 0 4304 0 1 4080
box -16 -6 32 210
use FILL  FILL_5323
timestamp 1018054153
transform 1 0 4320 0 1 4080
box -16 -6 32 210
use FILL  FILL_5325
timestamp 1018054153
transform 1 0 4336 0 1 4080
box -16 -6 32 210
use FILL  FILL_5327
timestamp 1018054153
transform 1 0 4352 0 1 4080
box -16 -6 32 210
use FILL  FILL_5329
timestamp 1018054153
transform 1 0 4368 0 1 4080
box -16 -6 32 210
use FILL  FILL_5331
timestamp 1018054153
transform 1 0 4384 0 1 4080
box -16 -6 32 210
use FILL  FILL_5333
timestamp 1018054153
transform 1 0 4400 0 1 4080
box -16 -6 32 210
use FILL  FILL_5335
timestamp 1018054153
transform 1 0 4416 0 1 4080
box -16 -6 32 210
use FILL  FILL_5337
timestamp 1018054153
transform 1 0 4432 0 1 4080
box -16 -6 32 210
use FILL  FILL_5339
timestamp 1018054153
transform 1 0 4448 0 1 4080
box -16 -6 32 210
use FILL  FILL_5341
timestamp 1018054153
transform 1 0 4464 0 1 4080
box -16 -6 32 210
use FILL  FILL_5343
timestamp 1018054153
transform 1 0 4480 0 1 4080
box -16 -6 32 210
use FILL  FILL_5345
timestamp 1018054153
transform 1 0 4496 0 1 4080
box -16 -6 32 210
use FILL  FILL_5347
timestamp 1018054153
transform 1 0 4512 0 1 4080
box -16 -6 32 210
use FILL  FILL_5349
timestamp 1018054153
transform 1 0 4528 0 1 4080
box -16 -6 32 210
use FILL  FILL_5351
timestamp 1018054153
transform 1 0 4544 0 1 4080
box -16 -6 32 210
use FILL  FILL_5353
timestamp 1018054153
transform 1 0 4560 0 1 4080
box -16 -6 32 210
use FILL  FILL_5355
timestamp 1018054153
transform 1 0 4576 0 1 4080
box -16 -6 32 210
use FILL  FILL_5357
timestamp 1018054153
transform 1 0 4592 0 1 4080
box -16 -6 32 210
use FILL  FILL_5359
timestamp 1018054153
transform 1 0 4608 0 1 4080
box -16 -6 32 210
use FILL  FILL_5361
timestamp 1018054153
transform 1 0 4624 0 1 4080
box -16 -6 32 210
use FILL  FILL_5363
timestamp 1018054153
transform 1 0 4640 0 1 4080
box -16 -6 32 210
use FILL  FILL_5365
timestamp 1018054153
transform 1 0 4656 0 1 4080
box -16 -6 32 210
use FILL  FILL_5367
timestamp 1018054153
transform 1 0 4672 0 1 4080
box -16 -6 32 210
use FILL  FILL_5369
timestamp 1018054153
transform 1 0 4688 0 1 4080
box -16 -6 32 210
use FILL  FILL_5371
timestamp 1018054153
transform 1 0 4704 0 1 4080
box -16 -6 32 210
use FILL  FILL_5373
timestamp 1018054153
transform 1 0 4720 0 1 4080
box -16 -6 32 210
use FILL  FILL_5375
timestamp 1018054153
transform 1 0 4736 0 1 4080
box -16 -6 32 210
use FILL  FILL_5377
timestamp 1018054153
transform 1 0 4752 0 1 4080
box -16 -6 32 210
use FILL  FILL_5379
timestamp 1018054153
transform 1 0 4768 0 1 4080
box -16 -6 32 210
use FILL  FILL_5381
timestamp 1018054153
transform 1 0 4784 0 1 4080
box -16 -6 32 210
use FILL  FILL_5383
timestamp 1018054153
transform 1 0 4800 0 1 4080
box -16 -6 32 210
use FILL  FILL_5385
timestamp 1018054153
transform 1 0 4816 0 1 4080
box -16 -6 32 210
use FILL  FILL_5387
timestamp 1018054153
transform 1 0 4832 0 1 4080
box -16 -6 32 210
use FILL  FILL_5389
timestamp 1018054153
transform 1 0 4848 0 1 4080
box -16 -6 32 210
use FILL  FILL_5391
timestamp 1018054153
transform 1 0 4864 0 1 4080
box -16 -6 32 210
use FILL  FILL_5393
timestamp 1018054153
transform 1 0 4880 0 1 4080
box -16 -6 32 210
use FILL  FILL_5395
timestamp 1018054153
transform 1 0 4896 0 1 4080
box -16 -6 32 210
use FILL  FILL_5397
timestamp 1018054153
transform 1 0 4912 0 1 4080
box -16 -6 32 210
use FILL  FILL_5399
timestamp 1018054153
transform 1 0 4928 0 1 4080
box -16 -6 32 210
use FILL  FILL_5401
timestamp 1018054153
transform 1 0 4944 0 1 4080
box -16 -6 32 210
use FILL  FILL_5403
timestamp 1018054153
transform 1 0 4960 0 1 4080
box -16 -6 32 210
use FILL  FILL_5405
timestamp 1018054153
transform 1 0 4976 0 1 4080
box -16 -6 32 210
use FILL  FILL_5407
timestamp 1018054153
transform 1 0 4992 0 1 4080
box -16 -6 32 210
use FILL  FILL_5409
timestamp 1018054153
transform 1 0 5008 0 1 4080
box -16 -6 32 210
use FILL  FILL_5411
timestamp 1018054153
transform 1 0 5024 0 1 4080
box -16 -6 32 210
use FILL  FILL_5413
timestamp 1018054153
transform 1 0 5040 0 1 4080
box -16 -6 32 210
use FILL  FILL_5414
timestamp 1018054153
transform 1 0 5056 0 1 4080
box -16 -6 32 210
use FILL  FILL_5415
timestamp 1018054153
transform 1 0 5072 0 1 4080
box -16 -6 32 210
use FILL  FILL_5416
timestamp 1018054153
transform 1 0 5088 0 1 4080
box -16 -6 32 210
use FILL  FILL_5417
timestamp 1018054153
transform 1 0 5104 0 1 4080
box -16 -6 32 210
use FILL  FILL_5418
timestamp 1018054153
transform 1 0 5120 0 1 4080
box -16 -6 32 210
use FILL  FILL_5419
timestamp 1018054153
transform 1 0 5136 0 1 4080
box -16 -6 32 210
use FILL  FILL_5420
timestamp 1018054153
transform 1 0 5152 0 1 4080
box -16 -6 32 210
use FILL  FILL_5421
timestamp 1018054153
transform 1 0 5168 0 1 4080
box -16 -6 32 210
use FILL  FILL_5422
timestamp 1018054153
transform 1 0 5184 0 1 4080
box -16 -6 32 210
use FILL  FILL_5423
timestamp 1018054153
transform 1 0 5200 0 1 4080
box -16 -6 32 210
use FILL  FILL_5424
timestamp 1018054153
transform 1 0 5216 0 1 4080
box -16 -6 32 210
use FILL  FILL_5425
timestamp 1018054153
transform 1 0 5232 0 1 4080
box -16 -6 32 210
use FILL  FILL_5426
timestamp 1018054153
transform 1 0 5248 0 1 4080
box -16 -6 32 210
use FILL  FILL_5427
timestamp 1018054153
transform 1 0 5264 0 1 4080
box -16 -6 32 210
use FILL  FILL_5428
timestamp 1018054153
transform 1 0 5280 0 1 4080
box -16 -6 32 210
use FILL  FILL_5429
timestamp 1018054153
transform 1 0 5296 0 1 4080
box -16 -6 32 210
use FILL  FILL_5430
timestamp 1018054153
transform 1 0 5312 0 1 4080
box -16 -6 32 210
use FILL  FILL_5431
timestamp 1018054153
transform 1 0 5328 0 1 4080
box -16 -6 32 210
use FILL  FILL_5432
timestamp 1018054153
transform 1 0 5344 0 1 4080
box -16 -6 32 210
use FILL  FILL_5433
timestamp 1018054153
transform 1 0 5360 0 1 4080
box -16 -6 32 210
use FILL  FILL_5434
timestamp 1018054153
transform 1 0 5376 0 1 4080
box -16 -6 32 210
use M3_M2  M3_M2_111
timestamp 1542725905
transform 1 0 5528 0 1 4090
box -6 -6 6 6
use M3_M2  M3_M2_112
timestamp 1542725905
transform 1 0 5560 0 1 4090
box -6 -6 6 6
use DFFSR  DFFSR_4
timestamp 1071163401
transform 1 0 5392 0 1 4080
box -16 -6 368 210
use FILL  FILL_5435
timestamp 1018054153
transform 1 0 5744 0 1 4080
box -16 -6 32 210
use FILL  FILL_5459
timestamp 1018054153
transform 1 0 5760 0 1 4080
box -16 -6 32 210
use FILL  FILL_5461
timestamp 1018054153
transform 1 0 5776 0 1 4080
box -16 -6 32 210
use FILL  FILL_5463
timestamp 1018054153
transform 1 0 5792 0 1 4080
box -16 -6 32 210
use FILL  FILL_5465
timestamp 1018054153
transform 1 0 5808 0 1 4080
box -16 -6 32 210
use FILL  FILL_5466
timestamp 1018054153
transform 1 0 5824 0 1 4080
box -16 -6 32 210
use FILL  FILL_5467
timestamp 1018054153
transform 1 0 5840 0 1 4080
box -16 -6 32 210
use FILL  FILL_5468
timestamp 1018054153
transform 1 0 5856 0 1 4080
box -16 -6 32 210
use FILL  FILL_5469
timestamp 1018054153
transform 1 0 5872 0 1 4080
box -16 -6 32 210
use FILL  FILL_5470
timestamp 1018054153
transform 1 0 5888 0 1 4080
box -16 -6 32 210
use FILL  FILL_5471
timestamp 1018054153
transform 1 0 5904 0 1 4080
box -16 -6 32 210
use FILL  FILL_5472
timestamp 1018054153
transform 1 0 5920 0 1 4080
box -16 -6 32 210
use FILL  FILL_5473
timestamp 1018054153
transform 1 0 5936 0 1 4080
box -16 -6 32 210
use FILL  FILL_5474
timestamp 1018054153
transform 1 0 5952 0 1 4080
box -16 -6 32 210
use FILL  FILL_5475
timestamp 1018054153
transform 1 0 5968 0 1 4080
box -16 -6 32 210
use FILL  FILL_5476
timestamp 1018054153
transform 1 0 5984 0 1 4080
box -16 -6 32 210
use FILL  FILL_5477
timestamp 1018054153
transform 1 0 6000 0 1 4080
box -16 -6 32 210
use FILL  FILL_5478
timestamp 1018054153
transform 1 0 6016 0 1 4080
box -16 -6 32 210
use FILL  FILL_5479
timestamp 1018054153
transform 1 0 6032 0 1 4080
box -16 -6 32 210
use FILL  FILL_5480
timestamp 1018054153
transform 1 0 6048 0 1 4080
box -16 -6 32 210
use FILL  FILL_5481
timestamp 1018054153
transform 1 0 6064 0 1 4080
box -16 -6 32 210
use BUFX2  BUFX2_3
timestamp 1090542073
transform 1 0 6080 0 1 4080
box -10 -6 56 210
use FILL  FILL_5482
timestamp 1018054153
transform 1 0 6128 0 1 4080
box -16 -6 32 210
use FILL  FILL_5483
timestamp 1018054153
transform 1 0 6144 0 1 4080
box -16 -6 32 210
use FILL  FILL_5484
timestamp 1018054153
transform 1 0 6160 0 1 4080
box -16 -6 32 210
use FILL  FILL_5486
timestamp 1018054153
transform 1 0 6176 0 1 4080
box -16 -6 32 210
use FILL  FILL_5488
timestamp 1018054153
transform 1 0 6192 0 1 4080
box -16 -6 32 210
use FILL  FILL_5490
timestamp 1018054153
transform 1 0 6208 0 1 4080
box -16 -6 32 210
use FILL  FILL_5492
timestamp 1018054153
transform 1 0 6224 0 1 4080
box -16 -6 32 210
use FILL  FILL_5494
timestamp 1018054153
transform 1 0 6240 0 1 4080
box -16 -6 32 210
use FILL  FILL_5496
timestamp 1018054153
transform 1 0 6256 0 1 4080
box -16 -6 32 210
use FILL  FILL_5498
timestamp 1018054153
transform 1 0 6272 0 1 4080
box -16 -6 32 210
use FILL  FILL_5500
timestamp 1018054153
transform 1 0 6288 0 1 4080
box -16 -6 32 210
use FILL  FILL_5502
timestamp 1018054153
transform 1 0 6304 0 1 4080
box -16 -6 32 210
use FILL  FILL_5504
timestamp 1018054153
transform 1 0 6320 0 1 4080
box -16 -6 32 210
use FILL  FILL_5506
timestamp 1018054153
transform 1 0 6336 0 1 4080
box -16 -6 32 210
use FILL  FILL_5508
timestamp 1018054153
transform 1 0 6352 0 1 4080
box -16 -6 32 210
use FILL  FILL_5510
timestamp 1018054153
transform 1 0 6368 0 1 4080
box -16 -6 32 210
use FILL  FILL_5512
timestamp 1018054153
transform 1 0 6384 0 1 4080
box -16 -6 32 210
use FILL  FILL_5514
timestamp 1018054153
transform 1 0 6400 0 1 4080
box -16 -6 32 210
use FILL  FILL_5516
timestamp 1018054153
transform 1 0 6416 0 1 4080
box -16 -6 32 210
use FILL  FILL_5518
timestamp 1018054153
transform 1 0 6432 0 1 4080
box -16 -6 32 210
use FILL  FILL_5520
timestamp 1018054153
transform 1 0 6448 0 1 4080
box -16 -6 32 210
use FILL  FILL_5522
timestamp 1018054153
transform 1 0 6464 0 1 4080
box -16 -6 32 210
use FILL  FILL_5524
timestamp 1018054153
transform 1 0 6480 0 1 4080
box -16 -6 32 210
use FILL  FILL_5526
timestamp 1018054153
transform 1 0 6496 0 1 4080
box -16 -6 32 210
use FILL  FILL_5528
timestamp 1018054153
transform 1 0 6512 0 1 4080
box -16 -6 32 210
use FILL  FILL_5530
timestamp 1018054153
transform 1 0 6528 0 1 4080
box -16 -6 32 210
use FILL  FILL_5532
timestamp 1018054153
transform 1 0 6544 0 1 4080
box -16 -6 32 210
use FILL  FILL_5534
timestamp 1018054153
transform 1 0 6560 0 1 4080
box -16 -6 32 210
use FILL  FILL_5536
timestamp 1018054153
transform 1 0 6576 0 1 4080
box -16 -6 32 210
use FILL  FILL_5538
timestamp 1018054153
transform 1 0 6592 0 1 4080
box -16 -6 32 210
use FILL  FILL_5540
timestamp 1018054153
transform 1 0 6608 0 1 4080
box -16 -6 32 210
use FILL  FILL_5542
timestamp 1018054153
transform 1 0 6624 0 1 4080
box -16 -6 32 210
use FILL  FILL_5544
timestamp 1018054153
transform 1 0 6640 0 1 4080
box -16 -6 32 210
use FILL  FILL_5546
timestamp 1018054153
transform 1 0 6656 0 1 4080
box -16 -6 32 210
use FILL  FILL_5548
timestamp 1018054153
transform 1 0 6672 0 1 4080
box -16 -6 32 210
use FILL  FILL_5550
timestamp 1018054153
transform 1 0 6688 0 1 4080
box -16 -6 32 210
use FILL  FILL_5552
timestamp 1018054153
transform 1 0 6704 0 1 4080
box -16 -6 32 210
use FILL  FILL_5554
timestamp 1018054153
transform 1 0 6720 0 1 4080
box -16 -6 32 210
use FILL  FILL_5556
timestamp 1018054153
transform 1 0 6736 0 1 4080
box -16 -6 32 210
use FILL  FILL_5558
timestamp 1018054153
transform 1 0 6752 0 1 4080
box -16 -6 32 210
use FILL  FILL_5560
timestamp 1018054153
transform 1 0 6768 0 1 4080
box -16 -6 32 210
use FILL  FILL_5562
timestamp 1018054153
transform 1 0 6784 0 1 4080
box -16 -6 32 210
use FILL  FILL_5563
timestamp 1018054153
transform 1 0 6800 0 1 4080
box -16 -6 32 210
use FILL  FILL_5564
timestamp 1018054153
transform 1 0 6816 0 1 4080
box -16 -6 32 210
use FILL  FILL_5565
timestamp 1018054153
transform 1 0 6832 0 1 4080
box -16 -6 32 210
use FILL  FILL_5566
timestamp 1018054153
transform 1 0 6848 0 1 4080
box -16 -6 32 210
use FILL  FILL_5567
timestamp 1018054153
transform 1 0 6864 0 1 4080
box -16 -6 32 210
use FILL  FILL_5568
timestamp 1018054153
transform 1 0 6880 0 1 4080
box -16 -6 32 210
use FILL  FILL_5569
timestamp 1018054153
transform 1 0 6896 0 1 4080
box -16 -6 32 210
use FILL  FILL_5570
timestamp 1018054153
transform 1 0 6912 0 1 4080
box -16 -6 32 210
use FILL  FILL_5571
timestamp 1018054153
transform 1 0 6928 0 1 4080
box -16 -6 32 210
use FILL  FILL_5572
timestamp 1018054153
transform 1 0 6944 0 1 4080
box -16 -6 32 210
use FILL  FILL_5573
timestamp 1018054153
transform 1 0 6960 0 1 4080
box -16 -6 32 210
use FILL  FILL_5574
timestamp 1018054153
transform 1 0 6976 0 1 4080
box -16 -6 32 210
use FILL  FILL_5575
timestamp 1018054153
transform 1 0 6992 0 1 4080
box -16 -6 32 210
use FILL  FILL_5576
timestamp 1018054153
transform 1 0 7008 0 1 4080
box -16 -6 32 210
use FILL  FILL_5577
timestamp 1018054153
transform 1 0 7024 0 1 4080
box -16 -6 32 210
use FILL  FILL_5578
timestamp 1018054153
transform 1 0 7040 0 1 4080
box -16 -6 32 210
use FILL  FILL_5579
timestamp 1018054153
transform 1 0 7056 0 1 4080
box -16 -6 32 210
use FILL  FILL_5580
timestamp 1018054153
transform 1 0 7072 0 1 4080
box -16 -6 32 210
use FILL  FILL_5581
timestamp 1018054153
transform 1 0 7088 0 1 4080
box -16 -6 32 210
use FILL  FILL_5582
timestamp 1018054153
transform 1 0 7104 0 1 4080
box -16 -6 32 210
use FILL  FILL_5583
timestamp 1018054153
transform 1 0 7120 0 1 4080
box -16 -6 32 210
use FILL  FILL_5584
timestamp 1018054153
transform 1 0 7136 0 1 4080
box -16 -6 32 210
use FILL  FILL_5586
timestamp 1018054153
transform 1 0 7152 0 1 4080
box -16 -6 32 210
use FILL  FILL_5588
timestamp 1018054153
transform 1 0 7168 0 1 4080
box -16 -6 32 210
use FILL  FILL_5590
timestamp 1018054153
transform 1 0 7184 0 1 4080
box -16 -6 32 210
use FILL  FILL_5592
timestamp 1018054153
transform 1 0 7200 0 1 4080
box -16 -6 32 210
use FILL  FILL_5594
timestamp 1018054153
transform 1 0 7216 0 1 4080
box -16 -6 32 210
use FILL  FILL_5596
timestamp 1018054153
transform 1 0 7232 0 1 4080
box -16 -6 32 210
use FILL  FILL_5598
timestamp 1018054153
transform 1 0 7248 0 1 4080
box -16 -6 32 210
use FILL  FILL_5600
timestamp 1018054153
transform 1 0 7264 0 1 4080
box -16 -6 32 210
use FILL  FILL_5602
timestamp 1018054153
transform 1 0 7280 0 1 4080
box -16 -6 32 210
use FILL  FILL_5604
timestamp 1018054153
transform 1 0 7296 0 1 4080
box -16 -6 32 210
use FILL  FILL_5606
timestamp 1018054153
transform 1 0 7312 0 1 4080
box -16 -6 32 210
use FILL  FILL_5608
timestamp 1018054153
transform 1 0 7328 0 1 4080
box -16 -6 32 210
use FILL  FILL_5610
timestamp 1018054153
transform 1 0 7344 0 1 4080
box -16 -6 32 210
use FILL  FILL_5612
timestamp 1018054153
transform 1 0 7360 0 1 4080
box -16 -6 32 210
use FILL  FILL_5614
timestamp 1018054153
transform 1 0 7376 0 1 4080
box -16 -6 32 210
use FILL  FILL_5616
timestamp 1018054153
transform 1 0 7392 0 1 4080
box -16 -6 32 210
use FILL  FILL_5618
timestamp 1018054153
transform 1 0 7408 0 1 4080
box -16 -6 32 210
use FILL  FILL_5620
timestamp 1018054153
transform 1 0 7424 0 1 4080
box -16 -6 32 210
use FILL  FILL_5622
timestamp 1018054153
transform 1 0 7440 0 1 4080
box -16 -6 32 210
use FILL  FILL_5624
timestamp 1018054153
transform 1 0 7456 0 1 4080
box -16 -6 32 210
use FILL  FILL_5626
timestamp 1018054153
transform 1 0 7472 0 1 4080
box -16 -6 32 210
use FILL  FILL_5628
timestamp 1018054153
transform 1 0 7488 0 1 4080
box -16 -6 32 210
use FILL  FILL_5630
timestamp 1018054153
transform 1 0 7504 0 1 4080
box -16 -6 32 210
use FILL  FILL_5632
timestamp 1018054153
transform 1 0 7520 0 1 4080
box -16 -6 32 210
use FILL  FILL_5634
timestamp 1018054153
transform 1 0 7536 0 1 4080
box -16 -6 32 210
use FILL  FILL_5636
timestamp 1018054153
transform 1 0 7552 0 1 4080
box -16 -6 32 210
use FILL  FILL_5638
timestamp 1018054153
transform 1 0 7568 0 1 4080
box -16 -6 32 210
use FILL  FILL_5640
timestamp 1018054153
transform 1 0 7584 0 1 4080
box -16 -6 32 210
use FILL  FILL_5642
timestamp 1018054153
transform 1 0 7600 0 1 4080
box -16 -6 32 210
use FILL  FILL_5644
timestamp 1018054153
transform 1 0 7616 0 1 4080
box -16 -6 32 210
use FILL  FILL_5646
timestamp 1018054153
transform 1 0 7632 0 1 4080
box -16 -6 32 210
use FILL  FILL_5648
timestamp 1018054153
transform 1 0 7648 0 1 4080
box -16 -6 32 210
use FILL  FILL_5650
timestamp 1018054153
transform 1 0 7664 0 1 4080
box -16 -6 32 210
use FILL  FILL_5652
timestamp 1018054153
transform 1 0 7680 0 1 4080
box -16 -6 32 210
use FILL  FILL_5654
timestamp 1018054153
transform 1 0 7696 0 1 4080
box -16 -6 32 210
use FILL  FILL_5656
timestamp 1018054153
transform 1 0 7712 0 1 4080
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_33
timestamp 1542725905
transform 1 0 7908 0 1 4080
box -48 -6 48 6
use M2_M1  M2_M1_261
timestamp 1542725905
transform 1 0 5208 0 1 4030
box -4 -4 4 4
use M2_M1  M2_M1_264
timestamp 1542725905
transform 1 0 5176 0 1 4010
box -4 -4 4 4
use M2_M1  M2_M1_267
timestamp 1542725905
transform 1 0 5112 0 1 3990
box -4 -4 4 4
use M2_M1  M2_M1_270
timestamp 1542725905
transform 1 0 5064 0 1 3970
box -4 -4 4 4
use M2_M1  M2_M1_273
timestamp 1542725905
transform 1 0 5384 0 1 3950
box -4 -4 4 4
use M3_M2  M3_M2_113
timestamp 1542725905
transform 1 0 5992 0 1 4070
box -6 -6 6 6
use M3_M2  M3_M2_114
timestamp 1542725905
transform 1 0 5944 0 1 4050
box -6 -6 6 6
use M2_M1  M2_M1_262
timestamp 1542725905
transform 1 0 5976 0 1 4030
box -4 -4 4 4
use M2_M1  M2_M1_265
timestamp 1542725905
transform 1 0 5944 0 1 4010
box -4 -4 4 4
use M2_M1  M2_M1_268
timestamp 1542725905
transform 1 0 5880 0 1 3990
box -4 -4 4 4
use M2_M1  M2_M1_271
timestamp 1542725905
transform 1 0 5832 0 1 3970
box -4 -4 4 4
use M3_M2  M3_M2_117
timestamp 1542725905
transform 1 0 5880 0 1 3970
box -6 -6 6 6
use M3_M2  M3_M2_118
timestamp 1542725905
transform 1 0 6072 0 1 3970
box -6 -6 6 6
use M2_M1  M2_M1_274
timestamp 1542725905
transform 1 0 6168 0 1 3950
box -4 -4 4 4
use M3_M2  M3_M2_115
timestamp 1542725905
transform 1 0 6408 0 1 4030
box -6 -6 6 6
use M3_M2  M3_M2_116
timestamp 1542725905
transform 1 0 6920 0 1 4030
box -6 -6 6 6
use M2_M1  M2_M1_263
timestamp 1542725905
transform 1 0 6952 0 1 4030
box -4 -4 4 4
use M2_M1  M2_M1_266
timestamp 1542725905
transform 1 0 6920 0 1 4010
box -4 -4 4 4
use M2_M1  M2_M1_269
timestamp 1542725905
transform 1 0 6856 0 1 3990
box -4 -4 4 4
use M2_M1  M2_M1_272
timestamp 1542725905
transform 1 0 6824 0 1 3970
box -4 -4 4 4
use M3_M2  M3_M2_119
timestamp 1542725905
transform 1 0 6856 0 1 3970
box -6 -6 6 6
use M2_M1  M2_M1_275
timestamp 1542725905
transform 1 0 7112 0 1 3950
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_34
timestamp 1542725905
transform 1 0 2212 0 1 3880
box -48 -6 48 6
use PADINC  PADINC_8
timestamp 1084294328
transform 0 -1 2000 1 0 3800
box -12 -6 606 2000
use M3_M2  M3_M2_120
timestamp 1542725905
transform 1 0 1998 0 1 3730
box -6 -6 6 6
use FILL  FILL_5068
timestamp 1018054153
transform 1 0 2272 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5070
timestamp 1018054153
transform 1 0 2288 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5072
timestamp 1018054153
transform 1 0 2304 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5074
timestamp 1018054153
transform 1 0 2320 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5076
timestamp 1018054153
transform 1 0 2336 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5078
timestamp 1018054153
transform 1 0 2352 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5080
timestamp 1018054153
transform 1 0 2368 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5082
timestamp 1018054153
transform 1 0 2384 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5084
timestamp 1018054153
transform 1 0 2400 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5086
timestamp 1018054153
transform 1 0 2416 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5088
timestamp 1018054153
transform 1 0 2432 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5090
timestamp 1018054153
transform 1 0 2448 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5092
timestamp 1018054153
transform 1 0 2464 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5094
timestamp 1018054153
transform 1 0 2480 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5096
timestamp 1018054153
transform 1 0 2496 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5098
timestamp 1018054153
transform 1 0 2512 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5100
timestamp 1018054153
transform 1 0 2528 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5102
timestamp 1018054153
transform 1 0 2544 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5104
timestamp 1018054153
transform 1 0 2560 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5106
timestamp 1018054153
transform 1 0 2576 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5108
timestamp 1018054153
transform 1 0 2592 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5110
timestamp 1018054153
transform 1 0 2608 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5112
timestamp 1018054153
transform 1 0 2624 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5114
timestamp 1018054153
transform 1 0 2640 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5116
timestamp 1018054153
transform 1 0 2656 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5118
timestamp 1018054153
transform 1 0 2672 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5120
timestamp 1018054153
transform 1 0 2688 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5122
timestamp 1018054153
transform 1 0 2704 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5124
timestamp 1018054153
transform 1 0 2720 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5126
timestamp 1018054153
transform 1 0 2736 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5128
timestamp 1018054153
transform 1 0 2752 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5130
timestamp 1018054153
transform 1 0 2768 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5132
timestamp 1018054153
transform 1 0 2784 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5134
timestamp 1018054153
transform 1 0 2800 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5136
timestamp 1018054153
transform 1 0 2816 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5138
timestamp 1018054153
transform 1 0 2832 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5140
timestamp 1018054153
transform 1 0 2848 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5142
timestamp 1018054153
transform 1 0 2864 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5144
timestamp 1018054153
transform 1 0 2880 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5146
timestamp 1018054153
transform 1 0 2896 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5148
timestamp 1018054153
transform 1 0 2912 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5150
timestamp 1018054153
transform 1 0 2928 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5152
timestamp 1018054153
transform 1 0 2944 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5154
timestamp 1018054153
transform 1 0 2960 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5156
timestamp 1018054153
transform 1 0 2976 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5158
timestamp 1018054153
transform 1 0 2992 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5160
timestamp 1018054153
transform 1 0 3008 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5162
timestamp 1018054153
transform 1 0 3024 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5164
timestamp 1018054153
transform 1 0 3040 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5166
timestamp 1018054153
transform 1 0 3056 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5168
timestamp 1018054153
transform 1 0 3072 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5170
timestamp 1018054153
transform 1 0 3088 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5172
timestamp 1018054153
transform 1 0 3104 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5174
timestamp 1018054153
transform 1 0 3120 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5176
timestamp 1018054153
transform 1 0 3136 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5178
timestamp 1018054153
transform 1 0 3152 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5180
timestamp 1018054153
transform 1 0 3168 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5182
timestamp 1018054153
transform 1 0 3184 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5184
timestamp 1018054153
transform 1 0 3200 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5186
timestamp 1018054153
transform 1 0 3216 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5188
timestamp 1018054153
transform 1 0 3232 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5190
timestamp 1018054153
transform 1 0 3248 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5192
timestamp 1018054153
transform 1 0 3264 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5194
timestamp 1018054153
transform 1 0 3280 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5196
timestamp 1018054153
transform 1 0 3296 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5198
timestamp 1018054153
transform 1 0 3312 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5200
timestamp 1018054153
transform 1 0 3328 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5202
timestamp 1018054153
transform 1 0 3344 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5204
timestamp 1018054153
transform 1 0 3360 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5206
timestamp 1018054153
transform 1 0 3376 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5208
timestamp 1018054153
transform 1 0 3392 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5210
timestamp 1018054153
transform 1 0 3408 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5212
timestamp 1018054153
transform 1 0 3424 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5214
timestamp 1018054153
transform 1 0 3440 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5216
timestamp 1018054153
transform 1 0 3456 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5218
timestamp 1018054153
transform 1 0 3472 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5220
timestamp 1018054153
transform 1 0 3488 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5222
timestamp 1018054153
transform 1 0 3504 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5224
timestamp 1018054153
transform 1 0 3520 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5226
timestamp 1018054153
transform 1 0 3536 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5228
timestamp 1018054153
transform 1 0 3552 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5230
timestamp 1018054153
transform 1 0 3568 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5232
timestamp 1018054153
transform 1 0 3584 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5234
timestamp 1018054153
transform 1 0 3600 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5236
timestamp 1018054153
transform 1 0 3616 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5238
timestamp 1018054153
transform 1 0 3632 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5240
timestamp 1018054153
transform 1 0 3648 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5242
timestamp 1018054153
transform 1 0 3664 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5244
timestamp 1018054153
transform 1 0 3680 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5246
timestamp 1018054153
transform 1 0 3696 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5248
timestamp 1018054153
transform 1 0 3712 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5250
timestamp 1018054153
transform 1 0 3728 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5252
timestamp 1018054153
transform 1 0 3744 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5254
timestamp 1018054153
transform 1 0 3760 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5256
timestamp 1018054153
transform 1 0 3776 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5258
timestamp 1018054153
transform 1 0 3792 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5260
timestamp 1018054153
transform 1 0 3808 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5262
timestamp 1018054153
transform 1 0 3824 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5264
timestamp 1018054153
transform 1 0 3840 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5266
timestamp 1018054153
transform 1 0 3856 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5268
timestamp 1018054153
transform 1 0 3872 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5270
timestamp 1018054153
transform 1 0 3888 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5272
timestamp 1018054153
transform 1 0 3904 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5274
timestamp 1018054153
transform 1 0 3920 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5276
timestamp 1018054153
transform 1 0 3936 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5278
timestamp 1018054153
transform 1 0 3952 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5280
timestamp 1018054153
transform 1 0 3968 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5282
timestamp 1018054153
transform 1 0 3984 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5284
timestamp 1018054153
transform 1 0 4000 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5286
timestamp 1018054153
transform 1 0 4016 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5288
timestamp 1018054153
transform 1 0 4032 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5290
timestamp 1018054153
transform 1 0 4048 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5292
timestamp 1018054153
transform 1 0 4064 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5294
timestamp 1018054153
transform 1 0 4080 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5296
timestamp 1018054153
transform 1 0 4096 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5298
timestamp 1018054153
transform 1 0 4112 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5300
timestamp 1018054153
transform 1 0 4128 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5302
timestamp 1018054153
transform 1 0 4144 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5304
timestamp 1018054153
transform 1 0 4160 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5306
timestamp 1018054153
transform 1 0 4176 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5308
timestamp 1018054153
transform 1 0 4192 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5310
timestamp 1018054153
transform 1 0 4208 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5312
timestamp 1018054153
transform 1 0 4224 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5314
timestamp 1018054153
transform 1 0 4240 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5316
timestamp 1018054153
transform 1 0 4256 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5318
timestamp 1018054153
transform 1 0 4272 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5320
timestamp 1018054153
transform 1 0 4288 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5322
timestamp 1018054153
transform 1 0 4304 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5324
timestamp 1018054153
transform 1 0 4320 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5326
timestamp 1018054153
transform 1 0 4336 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5328
timestamp 1018054153
transform 1 0 4352 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5330
timestamp 1018054153
transform 1 0 4368 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5332
timestamp 1018054153
transform 1 0 4384 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5334
timestamp 1018054153
transform 1 0 4400 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5336
timestamp 1018054153
transform 1 0 4416 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5338
timestamp 1018054153
transform 1 0 4432 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5340
timestamp 1018054153
transform 1 0 4448 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5342
timestamp 1018054153
transform 1 0 4464 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5344
timestamp 1018054153
transform 1 0 4480 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5346
timestamp 1018054153
transform 1 0 4496 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5348
timestamp 1018054153
transform 1 0 4512 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5350
timestamp 1018054153
transform 1 0 4528 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5352
timestamp 1018054153
transform 1 0 4544 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5354
timestamp 1018054153
transform 1 0 4560 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5356
timestamp 1018054153
transform 1 0 4576 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5358
timestamp 1018054153
transform 1 0 4592 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5360
timestamp 1018054153
transform 1 0 4608 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5362
timestamp 1018054153
transform 1 0 4624 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5364
timestamp 1018054153
transform 1 0 4640 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5366
timestamp 1018054153
transform 1 0 4656 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5368
timestamp 1018054153
transform 1 0 4672 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5370
timestamp 1018054153
transform 1 0 4688 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5372
timestamp 1018054153
transform 1 0 4704 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5374
timestamp 1018054153
transform 1 0 4720 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5376
timestamp 1018054153
transform 1 0 4736 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5378
timestamp 1018054153
transform 1 0 4752 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5380
timestamp 1018054153
transform 1 0 4768 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5382
timestamp 1018054153
transform 1 0 4784 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5384
timestamp 1018054153
transform 1 0 4800 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5386
timestamp 1018054153
transform 1 0 4816 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5388
timestamp 1018054153
transform 1 0 4832 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5390
timestamp 1018054153
transform 1 0 4848 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5392
timestamp 1018054153
transform 1 0 4864 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5394
timestamp 1018054153
transform 1 0 4880 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5396
timestamp 1018054153
transform 1 0 4896 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5398
timestamp 1018054153
transform 1 0 4912 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5400
timestamp 1018054153
transform 1 0 4928 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5402
timestamp 1018054153
transform 1 0 4944 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5404
timestamp 1018054153
transform 1 0 4960 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5406
timestamp 1018054153
transform 1 0 4976 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5408
timestamp 1018054153
transform 1 0 4992 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5410
timestamp 1018054153
transform 1 0 5008 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5412
timestamp 1018054153
transform 1 0 5024 0 -1 4080
box -16 -6 32 210
use M2_M1  M2_M1_276
timestamp 1542725905
transform 1 0 5064 0 1 3880
box -4 -4 4 4
use DFFSR  DFFSR_5
timestamp 1071163401
transform 1 0 5040 0 -1 4080
box -16 -6 368 210
use FILL  FILL_5436
timestamp 1018054153
transform 1 0 5392 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5437
timestamp 1018054153
transform 1 0 5408 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5438
timestamp 1018054153
transform 1 0 5424 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5439
timestamp 1018054153
transform 1 0 5440 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5440
timestamp 1018054153
transform 1 0 5456 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5441
timestamp 1018054153
transform 1 0 5472 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5442
timestamp 1018054153
transform 1 0 5488 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5443
timestamp 1018054153
transform 1 0 5504 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5444
timestamp 1018054153
transform 1 0 5520 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5445
timestamp 1018054153
transform 1 0 5536 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5446
timestamp 1018054153
transform 1 0 5552 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5447
timestamp 1018054153
transform 1 0 5568 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5448
timestamp 1018054153
transform 1 0 5584 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5449
timestamp 1018054153
transform 1 0 5600 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5450
timestamp 1018054153
transform 1 0 5616 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5451
timestamp 1018054153
transform 1 0 5632 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5452
timestamp 1018054153
transform 1 0 5648 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5453
timestamp 1018054153
transform 1 0 5664 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5454
timestamp 1018054153
transform 1 0 5680 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5455
timestamp 1018054153
transform 1 0 5696 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5456
timestamp 1018054153
transform 1 0 5712 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5457
timestamp 1018054153
transform 1 0 5728 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5458
timestamp 1018054153
transform 1 0 5744 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5460
timestamp 1018054153
transform 1 0 5760 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5462
timestamp 1018054153
transform 1 0 5776 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5464
timestamp 1018054153
transform 1 0 5792 0 -1 4080
box -16 -6 32 210
use M2_M1  M2_M1_277
timestamp 1542725905
transform 1 0 5832 0 1 3880
box -4 -4 4 4
use DFFSR  DFFSR_6
timestamp 1071163401
transform 1 0 5808 0 -1 4080
box -16 -6 368 210
use FILL  FILL_5485
timestamp 1018054153
transform 1 0 6160 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5487
timestamp 1018054153
transform 1 0 6176 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5489
timestamp 1018054153
transform 1 0 6192 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5491
timestamp 1018054153
transform 1 0 6208 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5493
timestamp 1018054153
transform 1 0 6224 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5495
timestamp 1018054153
transform 1 0 6240 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5497
timestamp 1018054153
transform 1 0 6256 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5499
timestamp 1018054153
transform 1 0 6272 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5501
timestamp 1018054153
transform 1 0 6288 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5503
timestamp 1018054153
transform 1 0 6304 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5505
timestamp 1018054153
transform 1 0 6320 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5507
timestamp 1018054153
transform 1 0 6336 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5509
timestamp 1018054153
transform 1 0 6352 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5511
timestamp 1018054153
transform 1 0 6368 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5513
timestamp 1018054153
transform 1 0 6384 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5515
timestamp 1018054153
transform 1 0 6400 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5517
timestamp 1018054153
transform 1 0 6416 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5519
timestamp 1018054153
transform 1 0 6432 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5521
timestamp 1018054153
transform 1 0 6448 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5523
timestamp 1018054153
transform 1 0 6464 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5525
timestamp 1018054153
transform 1 0 6480 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5527
timestamp 1018054153
transform 1 0 6496 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5529
timestamp 1018054153
transform 1 0 6512 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5531
timestamp 1018054153
transform 1 0 6528 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5533
timestamp 1018054153
transform 1 0 6544 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5535
timestamp 1018054153
transform 1 0 6560 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5537
timestamp 1018054153
transform 1 0 6576 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5539
timestamp 1018054153
transform 1 0 6592 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5541
timestamp 1018054153
transform 1 0 6608 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5543
timestamp 1018054153
transform 1 0 6624 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5545
timestamp 1018054153
transform 1 0 6640 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5547
timestamp 1018054153
transform 1 0 6656 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5549
timestamp 1018054153
transform 1 0 6672 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5551
timestamp 1018054153
transform 1 0 6688 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5553
timestamp 1018054153
transform 1 0 6704 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5555
timestamp 1018054153
transform 1 0 6720 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5557
timestamp 1018054153
transform 1 0 6736 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5559
timestamp 1018054153
transform 1 0 6752 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5561
timestamp 1018054153
transform 1 0 6768 0 -1 4080
box -16 -6 32 210
use M2_M1  M2_M1_278
timestamp 1542725905
transform 1 0 6824 0 1 3880
box -4 -4 4 4
use DFFSR  DFFSR_7
timestamp 1071163401
transform 1 0 6784 0 -1 4080
box -16 -6 368 210
use FILL  FILL_5585
timestamp 1018054153
transform 1 0 7136 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5587
timestamp 1018054153
transform 1 0 7152 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5589
timestamp 1018054153
transform 1 0 7168 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5591
timestamp 1018054153
transform 1 0 7184 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5593
timestamp 1018054153
transform 1 0 7200 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5595
timestamp 1018054153
transform 1 0 7216 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5597
timestamp 1018054153
transform 1 0 7232 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5599
timestamp 1018054153
transform 1 0 7248 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5601
timestamp 1018054153
transform 1 0 7264 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5603
timestamp 1018054153
transform 1 0 7280 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5605
timestamp 1018054153
transform 1 0 7296 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5607
timestamp 1018054153
transform 1 0 7312 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5609
timestamp 1018054153
transform 1 0 7328 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5611
timestamp 1018054153
transform 1 0 7344 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5613
timestamp 1018054153
transform 1 0 7360 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5615
timestamp 1018054153
transform 1 0 7376 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5617
timestamp 1018054153
transform 1 0 7392 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5619
timestamp 1018054153
transform 1 0 7408 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5621
timestamp 1018054153
transform 1 0 7424 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5623
timestamp 1018054153
transform 1 0 7440 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5625
timestamp 1018054153
transform 1 0 7456 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5627
timestamp 1018054153
transform 1 0 7472 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5629
timestamp 1018054153
transform 1 0 7488 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5631
timestamp 1018054153
transform 1 0 7504 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5633
timestamp 1018054153
transform 1 0 7520 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5635
timestamp 1018054153
transform 1 0 7536 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5637
timestamp 1018054153
transform 1 0 7552 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5639
timestamp 1018054153
transform 1 0 7568 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5641
timestamp 1018054153
transform 1 0 7584 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5643
timestamp 1018054153
transform 1 0 7600 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5645
timestamp 1018054153
transform 1 0 7616 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5647
timestamp 1018054153
transform 1 0 7632 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5649
timestamp 1018054153
transform 1 0 7648 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5651
timestamp 1018054153
transform 1 0 7664 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5653
timestamp 1018054153
transform 1 0 7680 0 -1 4080
box -16 -6 32 210
use FILL  FILL_5655
timestamp 1018054153
transform 1 0 7696 0 -1 4080
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_35
timestamp 1542725905
transform 1 0 7788 0 1 3880
box -48 -6 48 6
use FILL  FILL_5657
timestamp 1018054153
transform 1 0 7712 0 -1 4080
box -16 -6 32 210
use M3_M2  M3_M2_121
timestamp 1542725905
transform 1 0 3528 0 1 3730
box -6 -6 6 6
use M2_M1  M2_M1_279
timestamp 1542725905
transform 1 0 5384 0 1 3770
box -4 -4 4 4
use M2_M1  M2_M1_280
timestamp 1542725905
transform 1 0 5768 0 1 3770
box -4 -4 4 4
use M3_M2  M3_M2_122
timestamp 1542725905
transform 1 0 5768 0 1 3710
box -6 -6 6 6
use M2_M1  M2_M1_282
timestamp 1542725905
transform 1 0 6600 0 1 3750
box -4 -4 4 4
use M2_M1  M2_M1_281
timestamp 1542725905
transform 1 0 7112 0 1 3770
box -4 -4 4 4
use PADOUT  PADOUT_2
timestamp 1084294529
transform 0 1 8000 -1 0 4400
box -12 -6 606 2000
use M3_M2  M3_M2_123
timestamp 1542725905
transform 1 0 8002 0 1 3710
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_36
timestamp 1542725905
transform 1 0 2092 0 1 3680
box -48 -6 48 6
use FILL  FILL_5658
timestamp 1018054153
transform 1 0 2272 0 1 3680
box -16 -6 32 210
use FILL  FILL_5660
timestamp 1018054153
transform 1 0 2288 0 1 3680
box -16 -6 32 210
use FILL  FILL_5662
timestamp 1018054153
transform 1 0 2304 0 1 3680
box -16 -6 32 210
use FILL  FILL_5664
timestamp 1018054153
transform 1 0 2320 0 1 3680
box -16 -6 32 210
use FILL  FILL_5666
timestamp 1018054153
transform 1 0 2336 0 1 3680
box -16 -6 32 210
use FILL  FILL_5668
timestamp 1018054153
transform 1 0 2352 0 1 3680
box -16 -6 32 210
use FILL  FILL_5670
timestamp 1018054153
transform 1 0 2368 0 1 3680
box -16 -6 32 210
use FILL  FILL_5672
timestamp 1018054153
transform 1 0 2384 0 1 3680
box -16 -6 32 210
use FILL  FILL_5674
timestamp 1018054153
transform 1 0 2400 0 1 3680
box -16 -6 32 210
use FILL  FILL_5676
timestamp 1018054153
transform 1 0 2416 0 1 3680
box -16 -6 32 210
use FILL  FILL_5678
timestamp 1018054153
transform 1 0 2432 0 1 3680
box -16 -6 32 210
use FILL  FILL_5680
timestamp 1018054153
transform 1 0 2448 0 1 3680
box -16 -6 32 210
use FILL  FILL_5682
timestamp 1018054153
transform 1 0 2464 0 1 3680
box -16 -6 32 210
use FILL  FILL_5684
timestamp 1018054153
transform 1 0 2480 0 1 3680
box -16 -6 32 210
use FILL  FILL_5686
timestamp 1018054153
transform 1 0 2496 0 1 3680
box -16 -6 32 210
use FILL  FILL_5688
timestamp 1018054153
transform 1 0 2512 0 1 3680
box -16 -6 32 210
use FILL  FILL_5690
timestamp 1018054153
transform 1 0 2528 0 1 3680
box -16 -6 32 210
use FILL  FILL_5692
timestamp 1018054153
transform 1 0 2544 0 1 3680
box -16 -6 32 210
use FILL  FILL_5694
timestamp 1018054153
transform 1 0 2560 0 1 3680
box -16 -6 32 210
use FILL  FILL_5696
timestamp 1018054153
transform 1 0 2576 0 1 3680
box -16 -6 32 210
use FILL  FILL_5698
timestamp 1018054153
transform 1 0 2592 0 1 3680
box -16 -6 32 210
use FILL  FILL_5700
timestamp 1018054153
transform 1 0 2608 0 1 3680
box -16 -6 32 210
use FILL  FILL_5702
timestamp 1018054153
transform 1 0 2624 0 1 3680
box -16 -6 32 210
use FILL  FILL_5704
timestamp 1018054153
transform 1 0 2640 0 1 3680
box -16 -6 32 210
use FILL  FILL_5706
timestamp 1018054153
transform 1 0 2656 0 1 3680
box -16 -6 32 210
use FILL  FILL_5708
timestamp 1018054153
transform 1 0 2672 0 1 3680
box -16 -6 32 210
use FILL  FILL_5710
timestamp 1018054153
transform 1 0 2688 0 1 3680
box -16 -6 32 210
use FILL  FILL_5712
timestamp 1018054153
transform 1 0 2704 0 1 3680
box -16 -6 32 210
use FILL  FILL_5714
timestamp 1018054153
transform 1 0 2720 0 1 3680
box -16 -6 32 210
use FILL  FILL_5716
timestamp 1018054153
transform 1 0 2736 0 1 3680
box -16 -6 32 210
use FILL  FILL_5718
timestamp 1018054153
transform 1 0 2752 0 1 3680
box -16 -6 32 210
use FILL  FILL_5720
timestamp 1018054153
transform 1 0 2768 0 1 3680
box -16 -6 32 210
use FILL  FILL_5722
timestamp 1018054153
transform 1 0 2784 0 1 3680
box -16 -6 32 210
use FILL  FILL_5724
timestamp 1018054153
transform 1 0 2800 0 1 3680
box -16 -6 32 210
use FILL  FILL_5726
timestamp 1018054153
transform 1 0 2816 0 1 3680
box -16 -6 32 210
use FILL  FILL_5728
timestamp 1018054153
transform 1 0 2832 0 1 3680
box -16 -6 32 210
use FILL  FILL_5730
timestamp 1018054153
transform 1 0 2848 0 1 3680
box -16 -6 32 210
use FILL  FILL_5732
timestamp 1018054153
transform 1 0 2864 0 1 3680
box -16 -6 32 210
use FILL  FILL_5734
timestamp 1018054153
transform 1 0 2880 0 1 3680
box -16 -6 32 210
use FILL  FILL_5736
timestamp 1018054153
transform 1 0 2896 0 1 3680
box -16 -6 32 210
use FILL  FILL_5738
timestamp 1018054153
transform 1 0 2912 0 1 3680
box -16 -6 32 210
use FILL  FILL_5740
timestamp 1018054153
transform 1 0 2928 0 1 3680
box -16 -6 32 210
use FILL  FILL_5742
timestamp 1018054153
transform 1 0 2944 0 1 3680
box -16 -6 32 210
use FILL  FILL_5744
timestamp 1018054153
transform 1 0 2960 0 1 3680
box -16 -6 32 210
use FILL  FILL_5746
timestamp 1018054153
transform 1 0 2976 0 1 3680
box -16 -6 32 210
use FILL  FILL_5748
timestamp 1018054153
transform 1 0 2992 0 1 3680
box -16 -6 32 210
use FILL  FILL_5750
timestamp 1018054153
transform 1 0 3008 0 1 3680
box -16 -6 32 210
use FILL  FILL_5752
timestamp 1018054153
transform 1 0 3024 0 1 3680
box -16 -6 32 210
use FILL  FILL_5754
timestamp 1018054153
transform 1 0 3040 0 1 3680
box -16 -6 32 210
use FILL  FILL_5756
timestamp 1018054153
transform 1 0 3056 0 1 3680
box -16 -6 32 210
use FILL  FILL_5758
timestamp 1018054153
transform 1 0 3072 0 1 3680
box -16 -6 32 210
use FILL  FILL_5760
timestamp 1018054153
transform 1 0 3088 0 1 3680
box -16 -6 32 210
use FILL  FILL_5762
timestamp 1018054153
transform 1 0 3104 0 1 3680
box -16 -6 32 210
use FILL  FILL_5764
timestamp 1018054153
transform 1 0 3120 0 1 3680
box -16 -6 32 210
use FILL  FILL_5766
timestamp 1018054153
transform 1 0 3136 0 1 3680
box -16 -6 32 210
use FILL  FILL_5768
timestamp 1018054153
transform 1 0 3152 0 1 3680
box -16 -6 32 210
use FILL  FILL_5770
timestamp 1018054153
transform 1 0 3168 0 1 3680
box -16 -6 32 210
use FILL  FILL_5772
timestamp 1018054153
transform 1 0 3184 0 1 3680
box -16 -6 32 210
use FILL  FILL_5774
timestamp 1018054153
transform 1 0 3200 0 1 3680
box -16 -6 32 210
use FILL  FILL_5776
timestamp 1018054153
transform 1 0 3216 0 1 3680
box -16 -6 32 210
use FILL  FILL_5778
timestamp 1018054153
transform 1 0 3232 0 1 3680
box -16 -6 32 210
use FILL  FILL_5780
timestamp 1018054153
transform 1 0 3248 0 1 3680
box -16 -6 32 210
use FILL  FILL_5782
timestamp 1018054153
transform 1 0 3264 0 1 3680
box -16 -6 32 210
use FILL  FILL_5784
timestamp 1018054153
transform 1 0 3280 0 1 3680
box -16 -6 32 210
use FILL  FILL_5786
timestamp 1018054153
transform 1 0 3296 0 1 3680
box -16 -6 32 210
use FILL  FILL_5788
timestamp 1018054153
transform 1 0 3312 0 1 3680
box -16 -6 32 210
use FILL  FILL_5790
timestamp 1018054153
transform 1 0 3328 0 1 3680
box -16 -6 32 210
use FILL  FILL_5792
timestamp 1018054153
transform 1 0 3344 0 1 3680
box -16 -6 32 210
use FILL  FILL_5794
timestamp 1018054153
transform 1 0 3360 0 1 3680
box -16 -6 32 210
use FILL  FILL_5796
timestamp 1018054153
transform 1 0 3376 0 1 3680
box -16 -6 32 210
use FILL  FILL_5798
timestamp 1018054153
transform 1 0 3392 0 1 3680
box -16 -6 32 210
use FILL  FILL_5800
timestamp 1018054153
transform 1 0 3408 0 1 3680
box -16 -6 32 210
use FILL  FILL_5802
timestamp 1018054153
transform 1 0 3424 0 1 3680
box -16 -6 32 210
use FILL  FILL_5804
timestamp 1018054153
transform 1 0 3440 0 1 3680
box -16 -6 32 210
use FILL  FILL_5806
timestamp 1018054153
transform 1 0 3456 0 1 3680
box -16 -6 32 210
use FILL  FILL_5808
timestamp 1018054153
transform 1 0 3472 0 1 3680
box -16 -6 32 210
use FILL  FILL_5810
timestamp 1018054153
transform 1 0 3488 0 1 3680
box -16 -6 32 210
use FILL  FILL_5812
timestamp 1018054153
transform 1 0 3504 0 1 3680
box -16 -6 32 210
use FILL  FILL_5814
timestamp 1018054153
transform 1 0 3520 0 1 3680
box -16 -6 32 210
use FILL  FILL_5816
timestamp 1018054153
transform 1 0 3536 0 1 3680
box -16 -6 32 210
use FILL  FILL_5818
timestamp 1018054153
transform 1 0 3552 0 1 3680
box -16 -6 32 210
use FILL  FILL_5820
timestamp 1018054153
transform 1 0 3568 0 1 3680
box -16 -6 32 210
use FILL  FILL_5822
timestamp 1018054153
transform 1 0 3584 0 1 3680
box -16 -6 32 210
use FILL  FILL_5824
timestamp 1018054153
transform 1 0 3600 0 1 3680
box -16 -6 32 210
use FILL  FILL_5826
timestamp 1018054153
transform 1 0 3616 0 1 3680
box -16 -6 32 210
use FILL  FILL_5828
timestamp 1018054153
transform 1 0 3632 0 1 3680
box -16 -6 32 210
use FILL  FILL_5830
timestamp 1018054153
transform 1 0 3648 0 1 3680
box -16 -6 32 210
use FILL  FILL_5832
timestamp 1018054153
transform 1 0 3664 0 1 3680
box -16 -6 32 210
use FILL  FILL_5834
timestamp 1018054153
transform 1 0 3680 0 1 3680
box -16 -6 32 210
use FILL  FILL_5836
timestamp 1018054153
transform 1 0 3696 0 1 3680
box -16 -6 32 210
use FILL  FILL_5838
timestamp 1018054153
transform 1 0 3712 0 1 3680
box -16 -6 32 210
use FILL  FILL_5840
timestamp 1018054153
transform 1 0 3728 0 1 3680
box -16 -6 32 210
use FILL  FILL_5842
timestamp 1018054153
transform 1 0 3744 0 1 3680
box -16 -6 32 210
use FILL  FILL_5844
timestamp 1018054153
transform 1 0 3760 0 1 3680
box -16 -6 32 210
use FILL  FILL_5846
timestamp 1018054153
transform 1 0 3776 0 1 3680
box -16 -6 32 210
use FILL  FILL_5848
timestamp 1018054153
transform 1 0 3792 0 1 3680
box -16 -6 32 210
use FILL  FILL_5850
timestamp 1018054153
transform 1 0 3808 0 1 3680
box -16 -6 32 210
use FILL  FILL_5852
timestamp 1018054153
transform 1 0 3824 0 1 3680
box -16 -6 32 210
use FILL  FILL_5854
timestamp 1018054153
transform 1 0 3840 0 1 3680
box -16 -6 32 210
use FILL  FILL_5856
timestamp 1018054153
transform 1 0 3856 0 1 3680
box -16 -6 32 210
use FILL  FILL_5858
timestamp 1018054153
transform 1 0 3872 0 1 3680
box -16 -6 32 210
use FILL  FILL_5860
timestamp 1018054153
transform 1 0 3888 0 1 3680
box -16 -6 32 210
use FILL  FILL_5862
timestamp 1018054153
transform 1 0 3904 0 1 3680
box -16 -6 32 210
use FILL  FILL_5864
timestamp 1018054153
transform 1 0 3920 0 1 3680
box -16 -6 32 210
use FILL  FILL_5866
timestamp 1018054153
transform 1 0 3936 0 1 3680
box -16 -6 32 210
use FILL  FILL_5868
timestamp 1018054153
transform 1 0 3952 0 1 3680
box -16 -6 32 210
use FILL  FILL_5870
timestamp 1018054153
transform 1 0 3968 0 1 3680
box -16 -6 32 210
use FILL  FILL_5872
timestamp 1018054153
transform 1 0 3984 0 1 3680
box -16 -6 32 210
use FILL  FILL_5874
timestamp 1018054153
transform 1 0 4000 0 1 3680
box -16 -6 32 210
use FILL  FILL_5876
timestamp 1018054153
transform 1 0 4016 0 1 3680
box -16 -6 32 210
use FILL  FILL_5878
timestamp 1018054153
transform 1 0 4032 0 1 3680
box -16 -6 32 210
use FILL  FILL_5880
timestamp 1018054153
transform 1 0 4048 0 1 3680
box -16 -6 32 210
use FILL  FILL_5882
timestamp 1018054153
transform 1 0 4064 0 1 3680
box -16 -6 32 210
use FILL  FILL_5884
timestamp 1018054153
transform 1 0 4080 0 1 3680
box -16 -6 32 210
use FILL  FILL_5886
timestamp 1018054153
transform 1 0 4096 0 1 3680
box -16 -6 32 210
use FILL  FILL_5888
timestamp 1018054153
transform 1 0 4112 0 1 3680
box -16 -6 32 210
use FILL  FILL_5890
timestamp 1018054153
transform 1 0 4128 0 1 3680
box -16 -6 32 210
use FILL  FILL_5892
timestamp 1018054153
transform 1 0 4144 0 1 3680
box -16 -6 32 210
use FILL  FILL_5894
timestamp 1018054153
transform 1 0 4160 0 1 3680
box -16 -6 32 210
use FILL  FILL_5896
timestamp 1018054153
transform 1 0 4176 0 1 3680
box -16 -6 32 210
use FILL  FILL_5898
timestamp 1018054153
transform 1 0 4192 0 1 3680
box -16 -6 32 210
use FILL  FILL_5900
timestamp 1018054153
transform 1 0 4208 0 1 3680
box -16 -6 32 210
use FILL  FILL_5902
timestamp 1018054153
transform 1 0 4224 0 1 3680
box -16 -6 32 210
use FILL  FILL_5904
timestamp 1018054153
transform 1 0 4240 0 1 3680
box -16 -6 32 210
use FILL  FILL_5906
timestamp 1018054153
transform 1 0 4256 0 1 3680
box -16 -6 32 210
use FILL  FILL_5908
timestamp 1018054153
transform 1 0 4272 0 1 3680
box -16 -6 32 210
use FILL  FILL_5910
timestamp 1018054153
transform 1 0 4288 0 1 3680
box -16 -6 32 210
use FILL  FILL_5912
timestamp 1018054153
transform 1 0 4304 0 1 3680
box -16 -6 32 210
use FILL  FILL_5914
timestamp 1018054153
transform 1 0 4320 0 1 3680
box -16 -6 32 210
use FILL  FILL_5916
timestamp 1018054153
transform 1 0 4336 0 1 3680
box -16 -6 32 210
use FILL  FILL_5918
timestamp 1018054153
transform 1 0 4352 0 1 3680
box -16 -6 32 210
use FILL  FILL_5920
timestamp 1018054153
transform 1 0 4368 0 1 3680
box -16 -6 32 210
use FILL  FILL_5922
timestamp 1018054153
transform 1 0 4384 0 1 3680
box -16 -6 32 210
use FILL  FILL_5924
timestamp 1018054153
transform 1 0 4400 0 1 3680
box -16 -6 32 210
use FILL  FILL_5926
timestamp 1018054153
transform 1 0 4416 0 1 3680
box -16 -6 32 210
use FILL  FILL_5928
timestamp 1018054153
transform 1 0 4432 0 1 3680
box -16 -6 32 210
use FILL  FILL_5930
timestamp 1018054153
transform 1 0 4448 0 1 3680
box -16 -6 32 210
use FILL  FILL_5932
timestamp 1018054153
transform 1 0 4464 0 1 3680
box -16 -6 32 210
use FILL  FILL_5934
timestamp 1018054153
transform 1 0 4480 0 1 3680
box -16 -6 32 210
use FILL  FILL_5936
timestamp 1018054153
transform 1 0 4496 0 1 3680
box -16 -6 32 210
use FILL  FILL_5938
timestamp 1018054153
transform 1 0 4512 0 1 3680
box -16 -6 32 210
use FILL  FILL_5940
timestamp 1018054153
transform 1 0 4528 0 1 3680
box -16 -6 32 210
use FILL  FILL_5942
timestamp 1018054153
transform 1 0 4544 0 1 3680
box -16 -6 32 210
use FILL  FILL_5944
timestamp 1018054153
transform 1 0 4560 0 1 3680
box -16 -6 32 210
use FILL  FILL_5946
timestamp 1018054153
transform 1 0 4576 0 1 3680
box -16 -6 32 210
use FILL  FILL_5948
timestamp 1018054153
transform 1 0 4592 0 1 3680
box -16 -6 32 210
use FILL  FILL_5950
timestamp 1018054153
transform 1 0 4608 0 1 3680
box -16 -6 32 210
use FILL  FILL_5952
timestamp 1018054153
transform 1 0 4624 0 1 3680
box -16 -6 32 210
use FILL  FILL_5954
timestamp 1018054153
transform 1 0 4640 0 1 3680
box -16 -6 32 210
use FILL  FILL_5956
timestamp 1018054153
transform 1 0 4656 0 1 3680
box -16 -6 32 210
use FILL  FILL_5958
timestamp 1018054153
transform 1 0 4672 0 1 3680
box -16 -6 32 210
use FILL  FILL_5960
timestamp 1018054153
transform 1 0 4688 0 1 3680
box -16 -6 32 210
use FILL  FILL_5962
timestamp 1018054153
transform 1 0 4704 0 1 3680
box -16 -6 32 210
use FILL  FILL_5964
timestamp 1018054153
transform 1 0 4720 0 1 3680
box -16 -6 32 210
use FILL  FILL_5966
timestamp 1018054153
transform 1 0 4736 0 1 3680
box -16 -6 32 210
use FILL  FILL_5968
timestamp 1018054153
transform 1 0 4752 0 1 3680
box -16 -6 32 210
use FILL  FILL_5970
timestamp 1018054153
transform 1 0 4768 0 1 3680
box -16 -6 32 210
use FILL  FILL_5972
timestamp 1018054153
transform 1 0 4784 0 1 3680
box -16 -6 32 210
use FILL  FILL_5974
timestamp 1018054153
transform 1 0 4800 0 1 3680
box -16 -6 32 210
use FILL  FILL_5976
timestamp 1018054153
transform 1 0 4816 0 1 3680
box -16 -6 32 210
use FILL  FILL_5978
timestamp 1018054153
transform 1 0 4832 0 1 3680
box -16 -6 32 210
use FILL  FILL_5980
timestamp 1018054153
transform 1 0 4848 0 1 3680
box -16 -6 32 210
use FILL  FILL_5982
timestamp 1018054153
transform 1 0 4864 0 1 3680
box -16 -6 32 210
use FILL  FILL_5984
timestamp 1018054153
transform 1 0 4880 0 1 3680
box -16 -6 32 210
use FILL  FILL_5986
timestamp 1018054153
transform 1 0 4896 0 1 3680
box -16 -6 32 210
use FILL  FILL_5988
timestamp 1018054153
transform 1 0 4912 0 1 3680
box -16 -6 32 210
use FILL  FILL_5990
timestamp 1018054153
transform 1 0 4928 0 1 3680
box -16 -6 32 210
use FILL  FILL_5992
timestamp 1018054153
transform 1 0 4944 0 1 3680
box -16 -6 32 210
use FILL  FILL_5994
timestamp 1018054153
transform 1 0 4960 0 1 3680
box -16 -6 32 210
use FILL  FILL_5996
timestamp 1018054153
transform 1 0 4976 0 1 3680
box -16 -6 32 210
use FILL  FILL_5998
timestamp 1018054153
transform 1 0 4992 0 1 3680
box -16 -6 32 210
use FILL  FILL_6000
timestamp 1018054153
transform 1 0 5008 0 1 3680
box -16 -6 32 210
use FILL  FILL_6002
timestamp 1018054153
transform 1 0 5024 0 1 3680
box -16 -6 32 210
use FILL  FILL_6004
timestamp 1018054153
transform 1 0 5040 0 1 3680
box -16 -6 32 210
use FILL  FILL_6006
timestamp 1018054153
transform 1 0 5056 0 1 3680
box -16 -6 32 210
use FILL  FILL_6008
timestamp 1018054153
transform 1 0 5072 0 1 3680
box -16 -6 32 210
use FILL  FILL_6010
timestamp 1018054153
transform 1 0 5088 0 1 3680
box -16 -6 32 210
use FILL  FILL_6012
timestamp 1018054153
transform 1 0 5104 0 1 3680
box -16 -6 32 210
use FILL  FILL_6014
timestamp 1018054153
transform 1 0 5120 0 1 3680
box -16 -6 32 210
use FILL  FILL_6016
timestamp 1018054153
transform 1 0 5136 0 1 3680
box -16 -6 32 210
use FILL  FILL_6018
timestamp 1018054153
transform 1 0 5152 0 1 3680
box -16 -6 32 210
use FILL  FILL_6020
timestamp 1018054153
transform 1 0 5168 0 1 3680
box -16 -6 32 210
use FILL  FILL_6022
timestamp 1018054153
transform 1 0 5184 0 1 3680
box -16 -6 32 210
use FILL  FILL_6024
timestamp 1018054153
transform 1 0 5200 0 1 3680
box -16 -6 32 210
use FILL  FILL_6026
timestamp 1018054153
transform 1 0 5216 0 1 3680
box -16 -6 32 210
use FILL  FILL_6028
timestamp 1018054153
transform 1 0 5232 0 1 3680
box -16 -6 32 210
use FILL  FILL_6030
timestamp 1018054153
transform 1 0 5248 0 1 3680
box -16 -6 32 210
use FILL  FILL_6032
timestamp 1018054153
transform 1 0 5264 0 1 3680
box -16 -6 32 210
use FILL  FILL_6034
timestamp 1018054153
transform 1 0 5280 0 1 3680
box -16 -6 32 210
use FILL  FILL_6036
timestamp 1018054153
transform 1 0 5296 0 1 3680
box -16 -6 32 210
use FILL  FILL_6038
timestamp 1018054153
transform 1 0 5312 0 1 3680
box -16 -6 32 210
use FILL  FILL_6040
timestamp 1018054153
transform 1 0 5328 0 1 3680
box -16 -6 32 210
use FILL  FILL_6042
timestamp 1018054153
transform 1 0 5344 0 1 3680
box -16 -6 32 210
use FILL  FILL_6044
timestamp 1018054153
transform 1 0 5360 0 1 3680
box -16 -6 32 210
use FILL  FILL_6046
timestamp 1018054153
transform 1 0 5376 0 1 3680
box -16 -6 32 210
use BUFX2  BUFX2_4
timestamp 1090542073
transform 1 0 5392 0 1 3680
box -10 -6 56 210
use FILL  FILL_6048
timestamp 1018054153
transform 1 0 5440 0 1 3680
box -16 -6 32 210
use FILL  FILL_6053
timestamp 1018054153
transform 1 0 5456 0 1 3680
box -16 -6 32 210
use FILL  FILL_6055
timestamp 1018054153
transform 1 0 5472 0 1 3680
box -16 -6 32 210
use FILL  FILL_6057
timestamp 1018054153
transform 1 0 5488 0 1 3680
box -16 -6 32 210
use FILL  FILL_6059
timestamp 1018054153
transform 1 0 5504 0 1 3680
box -16 -6 32 210
use FILL  FILL_6061
timestamp 1018054153
transform 1 0 5520 0 1 3680
box -16 -6 32 210
use FILL  FILL_6063
timestamp 1018054153
transform 1 0 5536 0 1 3680
box -16 -6 32 210
use FILL  FILL_6065
timestamp 1018054153
transform 1 0 5552 0 1 3680
box -16 -6 32 210
use FILL  FILL_6067
timestamp 1018054153
transform 1 0 5568 0 1 3680
box -16 -6 32 210
use FILL  FILL_6069
timestamp 1018054153
transform 1 0 5584 0 1 3680
box -16 -6 32 210
use FILL  FILL_6071
timestamp 1018054153
transform 1 0 5600 0 1 3680
box -16 -6 32 210
use FILL  FILL_6073
timestamp 1018054153
transform 1 0 5616 0 1 3680
box -16 -6 32 210
use FILL  FILL_6075
timestamp 1018054153
transform 1 0 5632 0 1 3680
box -16 -6 32 210
use FILL  FILL_6077
timestamp 1018054153
transform 1 0 5648 0 1 3680
box -16 -6 32 210
use FILL  FILL_6079
timestamp 1018054153
transform 1 0 5664 0 1 3680
box -16 -6 32 210
use FILL  FILL_6081
timestamp 1018054153
transform 1 0 5680 0 1 3680
box -16 -6 32 210
use FILL  FILL_6083
timestamp 1018054153
transform 1 0 5696 0 1 3680
box -16 -6 32 210
use FILL  FILL_6085
timestamp 1018054153
transform 1 0 5712 0 1 3680
box -16 -6 32 210
use FILL  FILL_6087
timestamp 1018054153
transform 1 0 5728 0 1 3680
box -16 -6 32 210
use FILL  FILL_6089
timestamp 1018054153
transform 1 0 5744 0 1 3680
box -16 -6 32 210
use FILL  FILL_6091
timestamp 1018054153
transform 1 0 5760 0 1 3680
box -16 -6 32 210
use FILL  FILL_6093
timestamp 1018054153
transform 1 0 5776 0 1 3680
box -16 -6 32 210
use FILL  FILL_6095
timestamp 1018054153
transform 1 0 5792 0 1 3680
box -16 -6 32 210
use FILL  FILL_6097
timestamp 1018054153
transform 1 0 5808 0 1 3680
box -16 -6 32 210
use FILL  FILL_6099
timestamp 1018054153
transform 1 0 5824 0 1 3680
box -16 -6 32 210
use FILL  FILL_6101
timestamp 1018054153
transform 1 0 5840 0 1 3680
box -16 -6 32 210
use FILL  FILL_6103
timestamp 1018054153
transform 1 0 5856 0 1 3680
box -16 -6 32 210
use FILL  FILL_6105
timestamp 1018054153
transform 1 0 5872 0 1 3680
box -16 -6 32 210
use FILL  FILL_6107
timestamp 1018054153
transform 1 0 5888 0 1 3680
box -16 -6 32 210
use FILL  FILL_6109
timestamp 1018054153
transform 1 0 5904 0 1 3680
box -16 -6 32 210
use FILL  FILL_6111
timestamp 1018054153
transform 1 0 5920 0 1 3680
box -16 -6 32 210
use FILL  FILL_6113
timestamp 1018054153
transform 1 0 5936 0 1 3680
box -16 -6 32 210
use FILL  FILL_6114
timestamp 1018054153
transform 1 0 5952 0 1 3680
box -16 -6 32 210
use FILL  FILL_6115
timestamp 1018054153
transform 1 0 5968 0 1 3680
box -16 -6 32 210
use FILL  FILL_6116
timestamp 1018054153
transform 1 0 5984 0 1 3680
box -16 -6 32 210
use FILL  FILL_6117
timestamp 1018054153
transform 1 0 6000 0 1 3680
box -16 -6 32 210
use FILL  FILL_6120
timestamp 1018054153
transform 1 0 6016 0 1 3680
box -16 -6 32 210
use FILL  FILL_6122
timestamp 1018054153
transform 1 0 6032 0 1 3680
box -16 -6 32 210
use FILL  FILL_6124
timestamp 1018054153
transform 1 0 6048 0 1 3680
box -16 -6 32 210
use FILL  FILL_6126
timestamp 1018054153
transform 1 0 6064 0 1 3680
box -16 -6 32 210
use FILL  FILL_6128
timestamp 1018054153
transform 1 0 6080 0 1 3680
box -16 -6 32 210
use FILL  FILL_6130
timestamp 1018054153
transform 1 0 6096 0 1 3680
box -16 -6 32 210
use FILL  FILL_6132
timestamp 1018054153
transform 1 0 6112 0 1 3680
box -16 -6 32 210
use FILL  FILL_6134
timestamp 1018054153
transform 1 0 6128 0 1 3680
box -16 -6 32 210
use FILL  FILL_6136
timestamp 1018054153
transform 1 0 6144 0 1 3680
box -16 -6 32 210
use FILL  FILL_6138
timestamp 1018054153
transform 1 0 6160 0 1 3680
box -16 -6 32 210
use FILL  FILL_6140
timestamp 1018054153
transform 1 0 6176 0 1 3680
box -16 -6 32 210
use FILL  FILL_6142
timestamp 1018054153
transform 1 0 6192 0 1 3680
box -16 -6 32 210
use FILL  FILL_6144
timestamp 1018054153
transform 1 0 6208 0 1 3680
box -16 -6 32 210
use FILL  FILL_6146
timestamp 1018054153
transform 1 0 6224 0 1 3680
box -16 -6 32 210
use FILL  FILL_6148
timestamp 1018054153
transform 1 0 6240 0 1 3680
box -16 -6 32 210
use FILL  FILL_6150
timestamp 1018054153
transform 1 0 6256 0 1 3680
box -16 -6 32 210
use FILL  FILL_6152
timestamp 1018054153
transform 1 0 6272 0 1 3680
box -16 -6 32 210
use FILL  FILL_6154
timestamp 1018054153
transform 1 0 6288 0 1 3680
box -16 -6 32 210
use FILL  FILL_6156
timestamp 1018054153
transform 1 0 6304 0 1 3680
box -16 -6 32 210
use FILL  FILL_6158
timestamp 1018054153
transform 1 0 6320 0 1 3680
box -16 -6 32 210
use FILL  FILL_6160
timestamp 1018054153
transform 1 0 6336 0 1 3680
box -16 -6 32 210
use FILL  FILL_6162
timestamp 1018054153
transform 1 0 6352 0 1 3680
box -16 -6 32 210
use FILL  FILL_6164
timestamp 1018054153
transform 1 0 6368 0 1 3680
box -16 -6 32 210
use FILL  FILL_6166
timestamp 1018054153
transform 1 0 6384 0 1 3680
box -16 -6 32 210
use FILL  FILL_6168
timestamp 1018054153
transform 1 0 6400 0 1 3680
box -16 -6 32 210
use FILL  FILL_6170
timestamp 1018054153
transform 1 0 6416 0 1 3680
box -16 -6 32 210
use FILL  FILL_6172
timestamp 1018054153
transform 1 0 6432 0 1 3680
box -16 -6 32 210
use FILL  FILL_6174
timestamp 1018054153
transform 1 0 6448 0 1 3680
box -16 -6 32 210
use FILL  FILL_6176
timestamp 1018054153
transform 1 0 6464 0 1 3680
box -16 -6 32 210
use FILL  FILL_6178
timestamp 1018054153
transform 1 0 6480 0 1 3680
box -16 -6 32 210
use FILL  FILL_6180
timestamp 1018054153
transform 1 0 6496 0 1 3680
box -16 -6 32 210
use FILL  FILL_6182
timestamp 1018054153
transform 1 0 6512 0 1 3680
box -16 -6 32 210
use FILL  FILL_6184
timestamp 1018054153
transform 1 0 6528 0 1 3680
box -16 -6 32 210
use FILL  FILL_6186
timestamp 1018054153
transform 1 0 6544 0 1 3680
box -16 -6 32 210
use FILL  FILL_6188
timestamp 1018054153
transform 1 0 6560 0 1 3680
box -16 -6 32 210
use FILL  FILL_6190
timestamp 1018054153
transform 1 0 6576 0 1 3680
box -16 -6 32 210
use BUFX2  BUFX2_6
timestamp 1090542073
transform -1 0 6640 0 1 3680
box -10 -6 56 210
use FILL  FILL_6191
timestamp 1018054153
transform 1 0 6640 0 1 3680
box -16 -6 32 210
use FILL  FILL_6197
timestamp 1018054153
transform 1 0 6656 0 1 3680
box -16 -6 32 210
use FILL  FILL_6199
timestamp 1018054153
transform 1 0 6672 0 1 3680
box -16 -6 32 210
use FILL  FILL_6201
timestamp 1018054153
transform 1 0 6688 0 1 3680
box -16 -6 32 210
use FILL  FILL_6203
timestamp 1018054153
transform 1 0 6704 0 1 3680
box -16 -6 32 210
use FILL  FILL_6205
timestamp 1018054153
transform 1 0 6720 0 1 3680
box -16 -6 32 210
use FILL  FILL_6207
timestamp 1018054153
transform 1 0 6736 0 1 3680
box -16 -6 32 210
use FILL  FILL_6209
timestamp 1018054153
transform 1 0 6752 0 1 3680
box -16 -6 32 210
use FILL  FILL_6211
timestamp 1018054153
transform 1 0 6768 0 1 3680
box -16 -6 32 210
use FILL  FILL_6213
timestamp 1018054153
transform 1 0 6784 0 1 3680
box -16 -6 32 210
use FILL  FILL_6215
timestamp 1018054153
transform 1 0 6800 0 1 3680
box -16 -6 32 210
use FILL  FILL_6217
timestamp 1018054153
transform 1 0 6816 0 1 3680
box -16 -6 32 210
use FILL  FILL_6219
timestamp 1018054153
transform 1 0 6832 0 1 3680
box -16 -6 32 210
use FILL  FILL_6221
timestamp 1018054153
transform 1 0 6848 0 1 3680
box -16 -6 32 210
use FILL  FILL_6223
timestamp 1018054153
transform 1 0 6864 0 1 3680
box -16 -6 32 210
use FILL  FILL_6225
timestamp 1018054153
transform 1 0 6880 0 1 3680
box -16 -6 32 210
use FILL  FILL_6227
timestamp 1018054153
transform 1 0 6896 0 1 3680
box -16 -6 32 210
use FILL  FILL_6229
timestamp 1018054153
transform 1 0 6912 0 1 3680
box -16 -6 32 210
use FILL  FILL_6231
timestamp 1018054153
transform 1 0 6928 0 1 3680
box -16 -6 32 210
use FILL  FILL_6233
timestamp 1018054153
transform 1 0 6944 0 1 3680
box -16 -6 32 210
use FILL  FILL_6235
timestamp 1018054153
transform 1 0 6960 0 1 3680
box -16 -6 32 210
use FILL  FILL_6237
timestamp 1018054153
transform 1 0 6976 0 1 3680
box -16 -6 32 210
use FILL  FILL_6239
timestamp 1018054153
transform 1 0 6992 0 1 3680
box -16 -6 32 210
use FILL  FILL_6241
timestamp 1018054153
transform 1 0 7008 0 1 3680
box -16 -6 32 210
use FILL  FILL_6243
timestamp 1018054153
transform 1 0 7024 0 1 3680
box -16 -6 32 210
use FILL  FILL_6245
timestamp 1018054153
transform 1 0 7040 0 1 3680
box -16 -6 32 210
use FILL  FILL_6247
timestamp 1018054153
transform 1 0 7056 0 1 3680
box -16 -6 32 210
use FILL  FILL_6249
timestamp 1018054153
transform 1 0 7072 0 1 3680
box -16 -6 32 210
use FILL  FILL_6251
timestamp 1018054153
transform 1 0 7088 0 1 3680
box -16 -6 32 210
use FILL  FILL_6253
timestamp 1018054153
transform 1 0 7104 0 1 3680
box -16 -6 32 210
use FILL  FILL_6255
timestamp 1018054153
transform 1 0 7120 0 1 3680
box -16 -6 32 210
use FILL  FILL_6257
timestamp 1018054153
transform 1 0 7136 0 1 3680
box -16 -6 32 210
use FILL  FILL_6259
timestamp 1018054153
transform 1 0 7152 0 1 3680
box -16 -6 32 210
use FILL  FILL_6261
timestamp 1018054153
transform 1 0 7168 0 1 3680
box -16 -6 32 210
use FILL  FILL_6263
timestamp 1018054153
transform 1 0 7184 0 1 3680
box -16 -6 32 210
use FILL  FILL_6265
timestamp 1018054153
transform 1 0 7200 0 1 3680
box -16 -6 32 210
use FILL  FILL_6267
timestamp 1018054153
transform 1 0 7216 0 1 3680
box -16 -6 32 210
use FILL  FILL_6269
timestamp 1018054153
transform 1 0 7232 0 1 3680
box -16 -6 32 210
use FILL  FILL_6271
timestamp 1018054153
transform 1 0 7248 0 1 3680
box -16 -6 32 210
use FILL  FILL_6273
timestamp 1018054153
transform 1 0 7264 0 1 3680
box -16 -6 32 210
use FILL  FILL_6275
timestamp 1018054153
transform 1 0 7280 0 1 3680
box -16 -6 32 210
use FILL  FILL_6277
timestamp 1018054153
transform 1 0 7296 0 1 3680
box -16 -6 32 210
use FILL  FILL_6279
timestamp 1018054153
transform 1 0 7312 0 1 3680
box -16 -6 32 210
use FILL  FILL_6281
timestamp 1018054153
transform 1 0 7328 0 1 3680
box -16 -6 32 210
use FILL  FILL_6283
timestamp 1018054153
transform 1 0 7344 0 1 3680
box -16 -6 32 210
use FILL  FILL_6285
timestamp 1018054153
transform 1 0 7360 0 1 3680
box -16 -6 32 210
use FILL  FILL_6287
timestamp 1018054153
transform 1 0 7376 0 1 3680
box -16 -6 32 210
use FILL  FILL_6289
timestamp 1018054153
transform 1 0 7392 0 1 3680
box -16 -6 32 210
use FILL  FILL_6291
timestamp 1018054153
transform 1 0 7408 0 1 3680
box -16 -6 32 210
use FILL  FILL_6293
timestamp 1018054153
transform 1 0 7424 0 1 3680
box -16 -6 32 210
use FILL  FILL_6295
timestamp 1018054153
transform 1 0 7440 0 1 3680
box -16 -6 32 210
use FILL  FILL_6297
timestamp 1018054153
transform 1 0 7456 0 1 3680
box -16 -6 32 210
use FILL  FILL_6299
timestamp 1018054153
transform 1 0 7472 0 1 3680
box -16 -6 32 210
use FILL  FILL_6301
timestamp 1018054153
transform 1 0 7488 0 1 3680
box -16 -6 32 210
use FILL  FILL_6303
timestamp 1018054153
transform 1 0 7504 0 1 3680
box -16 -6 32 210
use FILL  FILL_6305
timestamp 1018054153
transform 1 0 7520 0 1 3680
box -16 -6 32 210
use FILL  FILL_6307
timestamp 1018054153
transform 1 0 7536 0 1 3680
box -16 -6 32 210
use FILL  FILL_6309
timestamp 1018054153
transform 1 0 7552 0 1 3680
box -16 -6 32 210
use FILL  FILL_6311
timestamp 1018054153
transform 1 0 7568 0 1 3680
box -16 -6 32 210
use FILL  FILL_6313
timestamp 1018054153
transform 1 0 7584 0 1 3680
box -16 -6 32 210
use FILL  FILL_6315
timestamp 1018054153
transform 1 0 7600 0 1 3680
box -16 -6 32 210
use FILL  FILL_6317
timestamp 1018054153
transform 1 0 7616 0 1 3680
box -16 -6 32 210
use FILL  FILL_6319
timestamp 1018054153
transform 1 0 7632 0 1 3680
box -16 -6 32 210
use FILL  FILL_6321
timestamp 1018054153
transform 1 0 7648 0 1 3680
box -16 -6 32 210
use FILL  FILL_6323
timestamp 1018054153
transform 1 0 7664 0 1 3680
box -16 -6 32 210
use FILL  FILL_6325
timestamp 1018054153
transform 1 0 7680 0 1 3680
box -16 -6 32 210
use FILL  FILL_6327
timestamp 1018054153
transform 1 0 7696 0 1 3680
box -16 -6 32 210
use FILL  FILL_6329
timestamp 1018054153
transform 1 0 7712 0 1 3680
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_37
timestamp 1542725905
transform 1 0 7908 0 1 3680
box -48 -6 48 6
use M2_M1  M2_M1_283
timestamp 1542725905
transform 1 0 5848 0 1 3610
box -4 -4 4 4
use M2_M1  M2_M1_284
timestamp 1542725905
transform 1 0 5944 0 1 3610
box -4 -4 4 4
use M2_M1  M2_M1_285
timestamp 1542725905
transform 1 0 6168 0 1 3590
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_38
timestamp 1542725905
transform 1 0 2212 0 1 3480
box -48 -6 48 6
use FILL  FILL_5659
timestamp 1018054153
transform 1 0 2272 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5661
timestamp 1018054153
transform 1 0 2288 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5663
timestamp 1018054153
transform 1 0 2304 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5665
timestamp 1018054153
transform 1 0 2320 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5667
timestamp 1018054153
transform 1 0 2336 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5669
timestamp 1018054153
transform 1 0 2352 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5671
timestamp 1018054153
transform 1 0 2368 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5673
timestamp 1018054153
transform 1 0 2384 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5675
timestamp 1018054153
transform 1 0 2400 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5677
timestamp 1018054153
transform 1 0 2416 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5679
timestamp 1018054153
transform 1 0 2432 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5681
timestamp 1018054153
transform 1 0 2448 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5683
timestamp 1018054153
transform 1 0 2464 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5685
timestamp 1018054153
transform 1 0 2480 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5687
timestamp 1018054153
transform 1 0 2496 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5689
timestamp 1018054153
transform 1 0 2512 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5691
timestamp 1018054153
transform 1 0 2528 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5693
timestamp 1018054153
transform 1 0 2544 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5695
timestamp 1018054153
transform 1 0 2560 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5697
timestamp 1018054153
transform 1 0 2576 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5699
timestamp 1018054153
transform 1 0 2592 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5701
timestamp 1018054153
transform 1 0 2608 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5703
timestamp 1018054153
transform 1 0 2624 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5705
timestamp 1018054153
transform 1 0 2640 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5707
timestamp 1018054153
transform 1 0 2656 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5709
timestamp 1018054153
transform 1 0 2672 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5711
timestamp 1018054153
transform 1 0 2688 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5713
timestamp 1018054153
transform 1 0 2704 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5715
timestamp 1018054153
transform 1 0 2720 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5717
timestamp 1018054153
transform 1 0 2736 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5719
timestamp 1018054153
transform 1 0 2752 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5721
timestamp 1018054153
transform 1 0 2768 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5723
timestamp 1018054153
transform 1 0 2784 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5725
timestamp 1018054153
transform 1 0 2800 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5727
timestamp 1018054153
transform 1 0 2816 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5729
timestamp 1018054153
transform 1 0 2832 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5731
timestamp 1018054153
transform 1 0 2848 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5733
timestamp 1018054153
transform 1 0 2864 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5735
timestamp 1018054153
transform 1 0 2880 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5737
timestamp 1018054153
transform 1 0 2896 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5739
timestamp 1018054153
transform 1 0 2912 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5741
timestamp 1018054153
transform 1 0 2928 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5743
timestamp 1018054153
transform 1 0 2944 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5745
timestamp 1018054153
transform 1 0 2960 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5747
timestamp 1018054153
transform 1 0 2976 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5749
timestamp 1018054153
transform 1 0 2992 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5751
timestamp 1018054153
transform 1 0 3008 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5753
timestamp 1018054153
transform 1 0 3024 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5755
timestamp 1018054153
transform 1 0 3040 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5757
timestamp 1018054153
transform 1 0 3056 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5759
timestamp 1018054153
transform 1 0 3072 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5761
timestamp 1018054153
transform 1 0 3088 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5763
timestamp 1018054153
transform 1 0 3104 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5765
timestamp 1018054153
transform 1 0 3120 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5767
timestamp 1018054153
transform 1 0 3136 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5769
timestamp 1018054153
transform 1 0 3152 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5771
timestamp 1018054153
transform 1 0 3168 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5773
timestamp 1018054153
transform 1 0 3184 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5775
timestamp 1018054153
transform 1 0 3200 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5777
timestamp 1018054153
transform 1 0 3216 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5779
timestamp 1018054153
transform 1 0 3232 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5781
timestamp 1018054153
transform 1 0 3248 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5783
timestamp 1018054153
transform 1 0 3264 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5785
timestamp 1018054153
transform 1 0 3280 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5787
timestamp 1018054153
transform 1 0 3296 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5789
timestamp 1018054153
transform 1 0 3312 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5791
timestamp 1018054153
transform 1 0 3328 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5793
timestamp 1018054153
transform 1 0 3344 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5795
timestamp 1018054153
transform 1 0 3360 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5797
timestamp 1018054153
transform 1 0 3376 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5799
timestamp 1018054153
transform 1 0 3392 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5801
timestamp 1018054153
transform 1 0 3408 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5803
timestamp 1018054153
transform 1 0 3424 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5805
timestamp 1018054153
transform 1 0 3440 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5807
timestamp 1018054153
transform 1 0 3456 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5809
timestamp 1018054153
transform 1 0 3472 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5811
timestamp 1018054153
transform 1 0 3488 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5813
timestamp 1018054153
transform 1 0 3504 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5815
timestamp 1018054153
transform 1 0 3520 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5817
timestamp 1018054153
transform 1 0 3536 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5819
timestamp 1018054153
transform 1 0 3552 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5821
timestamp 1018054153
transform 1 0 3568 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5823
timestamp 1018054153
transform 1 0 3584 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5825
timestamp 1018054153
transform 1 0 3600 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5827
timestamp 1018054153
transform 1 0 3616 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5829
timestamp 1018054153
transform 1 0 3632 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5831
timestamp 1018054153
transform 1 0 3648 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5833
timestamp 1018054153
transform 1 0 3664 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5835
timestamp 1018054153
transform 1 0 3680 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5837
timestamp 1018054153
transform 1 0 3696 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5839
timestamp 1018054153
transform 1 0 3712 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5841
timestamp 1018054153
transform 1 0 3728 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5843
timestamp 1018054153
transform 1 0 3744 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5845
timestamp 1018054153
transform 1 0 3760 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5847
timestamp 1018054153
transform 1 0 3776 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5849
timestamp 1018054153
transform 1 0 3792 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5851
timestamp 1018054153
transform 1 0 3808 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5853
timestamp 1018054153
transform 1 0 3824 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5855
timestamp 1018054153
transform 1 0 3840 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5857
timestamp 1018054153
transform 1 0 3856 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5859
timestamp 1018054153
transform 1 0 3872 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5861
timestamp 1018054153
transform 1 0 3888 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5863
timestamp 1018054153
transform 1 0 3904 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5865
timestamp 1018054153
transform 1 0 3920 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5867
timestamp 1018054153
transform 1 0 3936 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5869
timestamp 1018054153
transform 1 0 3952 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5871
timestamp 1018054153
transform 1 0 3968 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5873
timestamp 1018054153
transform 1 0 3984 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5875
timestamp 1018054153
transform 1 0 4000 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5877
timestamp 1018054153
transform 1 0 4016 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5879
timestamp 1018054153
transform 1 0 4032 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5881
timestamp 1018054153
transform 1 0 4048 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5883
timestamp 1018054153
transform 1 0 4064 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5885
timestamp 1018054153
transform 1 0 4080 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5887
timestamp 1018054153
transform 1 0 4096 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5889
timestamp 1018054153
transform 1 0 4112 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5891
timestamp 1018054153
transform 1 0 4128 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5893
timestamp 1018054153
transform 1 0 4144 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5895
timestamp 1018054153
transform 1 0 4160 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5897
timestamp 1018054153
transform 1 0 4176 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5899
timestamp 1018054153
transform 1 0 4192 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5901
timestamp 1018054153
transform 1 0 4208 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5903
timestamp 1018054153
transform 1 0 4224 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5905
timestamp 1018054153
transform 1 0 4240 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5907
timestamp 1018054153
transform 1 0 4256 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5909
timestamp 1018054153
transform 1 0 4272 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5911
timestamp 1018054153
transform 1 0 4288 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5913
timestamp 1018054153
transform 1 0 4304 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5915
timestamp 1018054153
transform 1 0 4320 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5917
timestamp 1018054153
transform 1 0 4336 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5919
timestamp 1018054153
transform 1 0 4352 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5921
timestamp 1018054153
transform 1 0 4368 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5923
timestamp 1018054153
transform 1 0 4384 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5925
timestamp 1018054153
transform 1 0 4400 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5927
timestamp 1018054153
transform 1 0 4416 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5929
timestamp 1018054153
transform 1 0 4432 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5931
timestamp 1018054153
transform 1 0 4448 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5933
timestamp 1018054153
transform 1 0 4464 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5935
timestamp 1018054153
transform 1 0 4480 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5937
timestamp 1018054153
transform 1 0 4496 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5939
timestamp 1018054153
transform 1 0 4512 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5941
timestamp 1018054153
transform 1 0 4528 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5943
timestamp 1018054153
transform 1 0 4544 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5945
timestamp 1018054153
transform 1 0 4560 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5947
timestamp 1018054153
transform 1 0 4576 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5949
timestamp 1018054153
transform 1 0 4592 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5951
timestamp 1018054153
transform 1 0 4608 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5953
timestamp 1018054153
transform 1 0 4624 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5955
timestamp 1018054153
transform 1 0 4640 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5957
timestamp 1018054153
transform 1 0 4656 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5959
timestamp 1018054153
transform 1 0 4672 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5961
timestamp 1018054153
transform 1 0 4688 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5963
timestamp 1018054153
transform 1 0 4704 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5965
timestamp 1018054153
transform 1 0 4720 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5967
timestamp 1018054153
transform 1 0 4736 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5969
timestamp 1018054153
transform 1 0 4752 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5971
timestamp 1018054153
transform 1 0 4768 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5973
timestamp 1018054153
transform 1 0 4784 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5975
timestamp 1018054153
transform 1 0 4800 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5977
timestamp 1018054153
transform 1 0 4816 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5979
timestamp 1018054153
transform 1 0 4832 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5981
timestamp 1018054153
transform 1 0 4848 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5983
timestamp 1018054153
transform 1 0 4864 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5985
timestamp 1018054153
transform 1 0 4880 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5987
timestamp 1018054153
transform 1 0 4896 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5989
timestamp 1018054153
transform 1 0 4912 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5991
timestamp 1018054153
transform 1 0 4928 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5993
timestamp 1018054153
transform 1 0 4944 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5995
timestamp 1018054153
transform 1 0 4960 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5997
timestamp 1018054153
transform 1 0 4976 0 -1 3680
box -16 -6 32 210
use FILL  FILL_5999
timestamp 1018054153
transform 1 0 4992 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6001
timestamp 1018054153
transform 1 0 5008 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6003
timestamp 1018054153
transform 1 0 5024 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6005
timestamp 1018054153
transform 1 0 5040 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6007
timestamp 1018054153
transform 1 0 5056 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6009
timestamp 1018054153
transform 1 0 5072 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6011
timestamp 1018054153
transform 1 0 5088 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6013
timestamp 1018054153
transform 1 0 5104 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6015
timestamp 1018054153
transform 1 0 5120 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6017
timestamp 1018054153
transform 1 0 5136 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6019
timestamp 1018054153
transform 1 0 5152 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6021
timestamp 1018054153
transform 1 0 5168 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6023
timestamp 1018054153
transform 1 0 5184 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6025
timestamp 1018054153
transform 1 0 5200 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6027
timestamp 1018054153
transform 1 0 5216 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6029
timestamp 1018054153
transform 1 0 5232 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6031
timestamp 1018054153
transform 1 0 5248 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6033
timestamp 1018054153
transform 1 0 5264 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6035
timestamp 1018054153
transform 1 0 5280 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6037
timestamp 1018054153
transform 1 0 5296 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6039
timestamp 1018054153
transform 1 0 5312 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6041
timestamp 1018054153
transform 1 0 5328 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6043
timestamp 1018054153
transform 1 0 5344 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6045
timestamp 1018054153
transform 1 0 5360 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6047
timestamp 1018054153
transform 1 0 5376 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6049
timestamp 1018054153
transform 1 0 5392 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6050
timestamp 1018054153
transform 1 0 5408 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6051
timestamp 1018054153
transform 1 0 5424 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6052
timestamp 1018054153
transform 1 0 5440 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6054
timestamp 1018054153
transform 1 0 5456 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6056
timestamp 1018054153
transform 1 0 5472 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6058
timestamp 1018054153
transform 1 0 5488 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6060
timestamp 1018054153
transform 1 0 5504 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6062
timestamp 1018054153
transform 1 0 5520 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6064
timestamp 1018054153
transform 1 0 5536 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6066
timestamp 1018054153
transform 1 0 5552 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6068
timestamp 1018054153
transform 1 0 5568 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6070
timestamp 1018054153
transform 1 0 5584 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6072
timestamp 1018054153
transform 1 0 5600 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6074
timestamp 1018054153
transform 1 0 5616 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6076
timestamp 1018054153
transform 1 0 5632 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6078
timestamp 1018054153
transform 1 0 5648 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6080
timestamp 1018054153
transform 1 0 5664 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6082
timestamp 1018054153
transform 1 0 5680 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6084
timestamp 1018054153
transform 1 0 5696 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6086
timestamp 1018054153
transform 1 0 5712 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6088
timestamp 1018054153
transform 1 0 5728 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6090
timestamp 1018054153
transform 1 0 5744 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6092
timestamp 1018054153
transform 1 0 5760 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6094
timestamp 1018054153
transform 1 0 5776 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6096
timestamp 1018054153
transform 1 0 5792 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6098
timestamp 1018054153
transform 1 0 5808 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6100
timestamp 1018054153
transform 1 0 5824 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6102
timestamp 1018054153
transform 1 0 5840 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6104
timestamp 1018054153
transform 1 0 5856 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6106
timestamp 1018054153
transform 1 0 5872 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6108
timestamp 1018054153
transform 1 0 5888 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6110
timestamp 1018054153
transform 1 0 5904 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6112
timestamp 1018054153
transform 1 0 5920 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6118
timestamp 1018054153
transform 1 0 5936 0 -1 3680
box -16 -6 32 210
use BUFX2  BUFX2_5
timestamp 1090542073
transform -1 0 6000 0 -1 3680
box -10 -6 56 210
use FILL  FILL_6119
timestamp 1018054153
transform 1 0 6000 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6121
timestamp 1018054153
transform 1 0 6016 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6123
timestamp 1018054153
transform 1 0 6032 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6125
timestamp 1018054153
transform 1 0 6048 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6127
timestamp 1018054153
transform 1 0 6064 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6129
timestamp 1018054153
transform 1 0 6080 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6131
timestamp 1018054153
transform 1 0 6096 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6133
timestamp 1018054153
transform 1 0 6112 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6135
timestamp 1018054153
transform 1 0 6128 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6137
timestamp 1018054153
transform 1 0 6144 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6139
timestamp 1018054153
transform 1 0 6160 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6141
timestamp 1018054153
transform 1 0 6176 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6143
timestamp 1018054153
transform 1 0 6192 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6145
timestamp 1018054153
transform 1 0 6208 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6147
timestamp 1018054153
transform 1 0 6224 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6149
timestamp 1018054153
transform 1 0 6240 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6151
timestamp 1018054153
transform 1 0 6256 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6153
timestamp 1018054153
transform 1 0 6272 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6155
timestamp 1018054153
transform 1 0 6288 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6157
timestamp 1018054153
transform 1 0 6304 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6159
timestamp 1018054153
transform 1 0 6320 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6161
timestamp 1018054153
transform 1 0 6336 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6163
timestamp 1018054153
transform 1 0 6352 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6165
timestamp 1018054153
transform 1 0 6368 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6167
timestamp 1018054153
transform 1 0 6384 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6169
timestamp 1018054153
transform 1 0 6400 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6171
timestamp 1018054153
transform 1 0 6416 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6173
timestamp 1018054153
transform 1 0 6432 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6175
timestamp 1018054153
transform 1 0 6448 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6177
timestamp 1018054153
transform 1 0 6464 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6179
timestamp 1018054153
transform 1 0 6480 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6181
timestamp 1018054153
transform 1 0 6496 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6183
timestamp 1018054153
transform 1 0 6512 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6185
timestamp 1018054153
transform 1 0 6528 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6187
timestamp 1018054153
transform 1 0 6544 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6189
timestamp 1018054153
transform 1 0 6560 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6192
timestamp 1018054153
transform 1 0 6576 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6193
timestamp 1018054153
transform 1 0 6592 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6194
timestamp 1018054153
transform 1 0 6608 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6195
timestamp 1018054153
transform 1 0 6624 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6196
timestamp 1018054153
transform 1 0 6640 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6198
timestamp 1018054153
transform 1 0 6656 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6200
timestamp 1018054153
transform 1 0 6672 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6202
timestamp 1018054153
transform 1 0 6688 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6204
timestamp 1018054153
transform 1 0 6704 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6206
timestamp 1018054153
transform 1 0 6720 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6208
timestamp 1018054153
transform 1 0 6736 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6210
timestamp 1018054153
transform 1 0 6752 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6212
timestamp 1018054153
transform 1 0 6768 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6214
timestamp 1018054153
transform 1 0 6784 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6216
timestamp 1018054153
transform 1 0 6800 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6218
timestamp 1018054153
transform 1 0 6816 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6220
timestamp 1018054153
transform 1 0 6832 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6222
timestamp 1018054153
transform 1 0 6848 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6224
timestamp 1018054153
transform 1 0 6864 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6226
timestamp 1018054153
transform 1 0 6880 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6228
timestamp 1018054153
transform 1 0 6896 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6230
timestamp 1018054153
transform 1 0 6912 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6232
timestamp 1018054153
transform 1 0 6928 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6234
timestamp 1018054153
transform 1 0 6944 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6236
timestamp 1018054153
transform 1 0 6960 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6238
timestamp 1018054153
transform 1 0 6976 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6240
timestamp 1018054153
transform 1 0 6992 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6242
timestamp 1018054153
transform 1 0 7008 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6244
timestamp 1018054153
transform 1 0 7024 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6246
timestamp 1018054153
transform 1 0 7040 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6248
timestamp 1018054153
transform 1 0 7056 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6250
timestamp 1018054153
transform 1 0 7072 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6252
timestamp 1018054153
transform 1 0 7088 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6254
timestamp 1018054153
transform 1 0 7104 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6256
timestamp 1018054153
transform 1 0 7120 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6258
timestamp 1018054153
transform 1 0 7136 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6260
timestamp 1018054153
transform 1 0 7152 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6262
timestamp 1018054153
transform 1 0 7168 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6264
timestamp 1018054153
transform 1 0 7184 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6266
timestamp 1018054153
transform 1 0 7200 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6268
timestamp 1018054153
transform 1 0 7216 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6270
timestamp 1018054153
transform 1 0 7232 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6272
timestamp 1018054153
transform 1 0 7248 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6274
timestamp 1018054153
transform 1 0 7264 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6276
timestamp 1018054153
transform 1 0 7280 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6278
timestamp 1018054153
transform 1 0 7296 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6280
timestamp 1018054153
transform 1 0 7312 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6282
timestamp 1018054153
transform 1 0 7328 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6284
timestamp 1018054153
transform 1 0 7344 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6286
timestamp 1018054153
transform 1 0 7360 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6288
timestamp 1018054153
transform 1 0 7376 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6290
timestamp 1018054153
transform 1 0 7392 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6292
timestamp 1018054153
transform 1 0 7408 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6294
timestamp 1018054153
transform 1 0 7424 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6296
timestamp 1018054153
transform 1 0 7440 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6298
timestamp 1018054153
transform 1 0 7456 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6300
timestamp 1018054153
transform 1 0 7472 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6302
timestamp 1018054153
transform 1 0 7488 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6304
timestamp 1018054153
transform 1 0 7504 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6306
timestamp 1018054153
transform 1 0 7520 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6308
timestamp 1018054153
transform 1 0 7536 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6310
timestamp 1018054153
transform 1 0 7552 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6312
timestamp 1018054153
transform 1 0 7568 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6314
timestamp 1018054153
transform 1 0 7584 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6316
timestamp 1018054153
transform 1 0 7600 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6318
timestamp 1018054153
transform 1 0 7616 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6320
timestamp 1018054153
transform 1 0 7632 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6322
timestamp 1018054153
transform 1 0 7648 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6324
timestamp 1018054153
transform 1 0 7664 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6326
timestamp 1018054153
transform 1 0 7680 0 -1 3680
box -16 -6 32 210
use FILL  FILL_6328
timestamp 1018054153
transform 1 0 7696 0 -1 3680
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_39
timestamp 1542725905
transform 1 0 7788 0 1 3480
box -48 -6 48 6
use FILL  FILL_6330
timestamp 1018054153
transform 1 0 7712 0 -1 3680
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_40
timestamp 1542725905
transform 1 0 2092 0 1 3280
box -48 -6 48 6
use FILL  FILL_6331
timestamp 1018054153
transform 1 0 2272 0 1 3280
box -16 -6 32 210
use FILL  FILL_6333
timestamp 1018054153
transform 1 0 2288 0 1 3280
box -16 -6 32 210
use FILL  FILL_6335
timestamp 1018054153
transform 1 0 2304 0 1 3280
box -16 -6 32 210
use FILL  FILL_6337
timestamp 1018054153
transform 1 0 2320 0 1 3280
box -16 -6 32 210
use FILL  FILL_6339
timestamp 1018054153
transform 1 0 2336 0 1 3280
box -16 -6 32 210
use FILL  FILL_6341
timestamp 1018054153
transform 1 0 2352 0 1 3280
box -16 -6 32 210
use FILL  FILL_6343
timestamp 1018054153
transform 1 0 2368 0 1 3280
box -16 -6 32 210
use FILL  FILL_6345
timestamp 1018054153
transform 1 0 2384 0 1 3280
box -16 -6 32 210
use FILL  FILL_6347
timestamp 1018054153
transform 1 0 2400 0 1 3280
box -16 -6 32 210
use FILL  FILL_6349
timestamp 1018054153
transform 1 0 2416 0 1 3280
box -16 -6 32 210
use FILL  FILL_6351
timestamp 1018054153
transform 1 0 2432 0 1 3280
box -16 -6 32 210
use FILL  FILL_6353
timestamp 1018054153
transform 1 0 2448 0 1 3280
box -16 -6 32 210
use FILL  FILL_6355
timestamp 1018054153
transform 1 0 2464 0 1 3280
box -16 -6 32 210
use FILL  FILL_6357
timestamp 1018054153
transform 1 0 2480 0 1 3280
box -16 -6 32 210
use FILL  FILL_6359
timestamp 1018054153
transform 1 0 2496 0 1 3280
box -16 -6 32 210
use FILL  FILL_6361
timestamp 1018054153
transform 1 0 2512 0 1 3280
box -16 -6 32 210
use FILL  FILL_6363
timestamp 1018054153
transform 1 0 2528 0 1 3280
box -16 -6 32 210
use FILL  FILL_6365
timestamp 1018054153
transform 1 0 2544 0 1 3280
box -16 -6 32 210
use FILL  FILL_6367
timestamp 1018054153
transform 1 0 2560 0 1 3280
box -16 -6 32 210
use FILL  FILL_6369
timestamp 1018054153
transform 1 0 2576 0 1 3280
box -16 -6 32 210
use FILL  FILL_6371
timestamp 1018054153
transform 1 0 2592 0 1 3280
box -16 -6 32 210
use FILL  FILL_6373
timestamp 1018054153
transform 1 0 2608 0 1 3280
box -16 -6 32 210
use FILL  FILL_6375
timestamp 1018054153
transform 1 0 2624 0 1 3280
box -16 -6 32 210
use FILL  FILL_6377
timestamp 1018054153
transform 1 0 2640 0 1 3280
box -16 -6 32 210
use FILL  FILL_6379
timestamp 1018054153
transform 1 0 2656 0 1 3280
box -16 -6 32 210
use FILL  FILL_6381
timestamp 1018054153
transform 1 0 2672 0 1 3280
box -16 -6 32 210
use FILL  FILL_6383
timestamp 1018054153
transform 1 0 2688 0 1 3280
box -16 -6 32 210
use FILL  FILL_6385
timestamp 1018054153
transform 1 0 2704 0 1 3280
box -16 -6 32 210
use FILL  FILL_6387
timestamp 1018054153
transform 1 0 2720 0 1 3280
box -16 -6 32 210
use FILL  FILL_6389
timestamp 1018054153
transform 1 0 2736 0 1 3280
box -16 -6 32 210
use FILL  FILL_6391
timestamp 1018054153
transform 1 0 2752 0 1 3280
box -16 -6 32 210
use FILL  FILL_6393
timestamp 1018054153
transform 1 0 2768 0 1 3280
box -16 -6 32 210
use FILL  FILL_6395
timestamp 1018054153
transform 1 0 2784 0 1 3280
box -16 -6 32 210
use FILL  FILL_6397
timestamp 1018054153
transform 1 0 2800 0 1 3280
box -16 -6 32 210
use FILL  FILL_6399
timestamp 1018054153
transform 1 0 2816 0 1 3280
box -16 -6 32 210
use FILL  FILL_6401
timestamp 1018054153
transform 1 0 2832 0 1 3280
box -16 -6 32 210
use FILL  FILL_6403
timestamp 1018054153
transform 1 0 2848 0 1 3280
box -16 -6 32 210
use FILL  FILL_6405
timestamp 1018054153
transform 1 0 2864 0 1 3280
box -16 -6 32 210
use FILL  FILL_6407
timestamp 1018054153
transform 1 0 2880 0 1 3280
box -16 -6 32 210
use FILL  FILL_6409
timestamp 1018054153
transform 1 0 2896 0 1 3280
box -16 -6 32 210
use FILL  FILL_6411
timestamp 1018054153
transform 1 0 2912 0 1 3280
box -16 -6 32 210
use FILL  FILL_6413
timestamp 1018054153
transform 1 0 2928 0 1 3280
box -16 -6 32 210
use FILL  FILL_6415
timestamp 1018054153
transform 1 0 2944 0 1 3280
box -16 -6 32 210
use FILL  FILL_6417
timestamp 1018054153
transform 1 0 2960 0 1 3280
box -16 -6 32 210
use FILL  FILL_6419
timestamp 1018054153
transform 1 0 2976 0 1 3280
box -16 -6 32 210
use FILL  FILL_6421
timestamp 1018054153
transform 1 0 2992 0 1 3280
box -16 -6 32 210
use FILL  FILL_6423
timestamp 1018054153
transform 1 0 3008 0 1 3280
box -16 -6 32 210
use FILL  FILL_6425
timestamp 1018054153
transform 1 0 3024 0 1 3280
box -16 -6 32 210
use FILL  FILL_6427
timestamp 1018054153
transform 1 0 3040 0 1 3280
box -16 -6 32 210
use FILL  FILL_6429
timestamp 1018054153
transform 1 0 3056 0 1 3280
box -16 -6 32 210
use FILL  FILL_6431
timestamp 1018054153
transform 1 0 3072 0 1 3280
box -16 -6 32 210
use FILL  FILL_6433
timestamp 1018054153
transform 1 0 3088 0 1 3280
box -16 -6 32 210
use FILL  FILL_6435
timestamp 1018054153
transform 1 0 3104 0 1 3280
box -16 -6 32 210
use FILL  FILL_6437
timestamp 1018054153
transform 1 0 3120 0 1 3280
box -16 -6 32 210
use FILL  FILL_6439
timestamp 1018054153
transform 1 0 3136 0 1 3280
box -16 -6 32 210
use FILL  FILL_6441
timestamp 1018054153
transform 1 0 3152 0 1 3280
box -16 -6 32 210
use FILL  FILL_6443
timestamp 1018054153
transform 1 0 3168 0 1 3280
box -16 -6 32 210
use FILL  FILL_6445
timestamp 1018054153
transform 1 0 3184 0 1 3280
box -16 -6 32 210
use FILL  FILL_6447
timestamp 1018054153
transform 1 0 3200 0 1 3280
box -16 -6 32 210
use FILL  FILL_6449
timestamp 1018054153
transform 1 0 3216 0 1 3280
box -16 -6 32 210
use FILL  FILL_6451
timestamp 1018054153
transform 1 0 3232 0 1 3280
box -16 -6 32 210
use FILL  FILL_6453
timestamp 1018054153
transform 1 0 3248 0 1 3280
box -16 -6 32 210
use FILL  FILL_6455
timestamp 1018054153
transform 1 0 3264 0 1 3280
box -16 -6 32 210
use FILL  FILL_6457
timestamp 1018054153
transform 1 0 3280 0 1 3280
box -16 -6 32 210
use FILL  FILL_6459
timestamp 1018054153
transform 1 0 3296 0 1 3280
box -16 -6 32 210
use FILL  FILL_6461
timestamp 1018054153
transform 1 0 3312 0 1 3280
box -16 -6 32 210
use FILL  FILL_6463
timestamp 1018054153
transform 1 0 3328 0 1 3280
box -16 -6 32 210
use FILL  FILL_6465
timestamp 1018054153
transform 1 0 3344 0 1 3280
box -16 -6 32 210
use FILL  FILL_6467
timestamp 1018054153
transform 1 0 3360 0 1 3280
box -16 -6 32 210
use FILL  FILL_6469
timestamp 1018054153
transform 1 0 3376 0 1 3280
box -16 -6 32 210
use FILL  FILL_6471
timestamp 1018054153
transform 1 0 3392 0 1 3280
box -16 -6 32 210
use FILL  FILL_6473
timestamp 1018054153
transform 1 0 3408 0 1 3280
box -16 -6 32 210
use FILL  FILL_6475
timestamp 1018054153
transform 1 0 3424 0 1 3280
box -16 -6 32 210
use FILL  FILL_6477
timestamp 1018054153
transform 1 0 3440 0 1 3280
box -16 -6 32 210
use FILL  FILL_6479
timestamp 1018054153
transform 1 0 3456 0 1 3280
box -16 -6 32 210
use FILL  FILL_6481
timestamp 1018054153
transform 1 0 3472 0 1 3280
box -16 -6 32 210
use FILL  FILL_6483
timestamp 1018054153
transform 1 0 3488 0 1 3280
box -16 -6 32 210
use FILL  FILL_6485
timestamp 1018054153
transform 1 0 3504 0 1 3280
box -16 -6 32 210
use FILL  FILL_6487
timestamp 1018054153
transform 1 0 3520 0 1 3280
box -16 -6 32 210
use FILL  FILL_6489
timestamp 1018054153
transform 1 0 3536 0 1 3280
box -16 -6 32 210
use FILL  FILL_6491
timestamp 1018054153
transform 1 0 3552 0 1 3280
box -16 -6 32 210
use FILL  FILL_6493
timestamp 1018054153
transform 1 0 3568 0 1 3280
box -16 -6 32 210
use FILL  FILL_6495
timestamp 1018054153
transform 1 0 3584 0 1 3280
box -16 -6 32 210
use FILL  FILL_6497
timestamp 1018054153
transform 1 0 3600 0 1 3280
box -16 -6 32 210
use FILL  FILL_6499
timestamp 1018054153
transform 1 0 3616 0 1 3280
box -16 -6 32 210
use FILL  FILL_6501
timestamp 1018054153
transform 1 0 3632 0 1 3280
box -16 -6 32 210
use FILL  FILL_6503
timestamp 1018054153
transform 1 0 3648 0 1 3280
box -16 -6 32 210
use FILL  FILL_6505
timestamp 1018054153
transform 1 0 3664 0 1 3280
box -16 -6 32 210
use FILL  FILL_6507
timestamp 1018054153
transform 1 0 3680 0 1 3280
box -16 -6 32 210
use FILL  FILL_6509
timestamp 1018054153
transform 1 0 3696 0 1 3280
box -16 -6 32 210
use FILL  FILL_6511
timestamp 1018054153
transform 1 0 3712 0 1 3280
box -16 -6 32 210
use FILL  FILL_6513
timestamp 1018054153
transform 1 0 3728 0 1 3280
box -16 -6 32 210
use FILL  FILL_6515
timestamp 1018054153
transform 1 0 3744 0 1 3280
box -16 -6 32 210
use FILL  FILL_6517
timestamp 1018054153
transform 1 0 3760 0 1 3280
box -16 -6 32 210
use FILL  FILL_6519
timestamp 1018054153
transform 1 0 3776 0 1 3280
box -16 -6 32 210
use FILL  FILL_6521
timestamp 1018054153
transform 1 0 3792 0 1 3280
box -16 -6 32 210
use FILL  FILL_6523
timestamp 1018054153
transform 1 0 3808 0 1 3280
box -16 -6 32 210
use FILL  FILL_6525
timestamp 1018054153
transform 1 0 3824 0 1 3280
box -16 -6 32 210
use FILL  FILL_6527
timestamp 1018054153
transform 1 0 3840 0 1 3280
box -16 -6 32 210
use FILL  FILL_6529
timestamp 1018054153
transform 1 0 3856 0 1 3280
box -16 -6 32 210
use FILL  FILL_6531
timestamp 1018054153
transform 1 0 3872 0 1 3280
box -16 -6 32 210
use FILL  FILL_6533
timestamp 1018054153
transform 1 0 3888 0 1 3280
box -16 -6 32 210
use FILL  FILL_6535
timestamp 1018054153
transform 1 0 3904 0 1 3280
box -16 -6 32 210
use FILL  FILL_6537
timestamp 1018054153
transform 1 0 3920 0 1 3280
box -16 -6 32 210
use FILL  FILL_6539
timestamp 1018054153
transform 1 0 3936 0 1 3280
box -16 -6 32 210
use FILL  FILL_6541
timestamp 1018054153
transform 1 0 3952 0 1 3280
box -16 -6 32 210
use FILL  FILL_6543
timestamp 1018054153
transform 1 0 3968 0 1 3280
box -16 -6 32 210
use FILL  FILL_6545
timestamp 1018054153
transform 1 0 3984 0 1 3280
box -16 -6 32 210
use FILL  FILL_6547
timestamp 1018054153
transform 1 0 4000 0 1 3280
box -16 -6 32 210
use FILL  FILL_6549
timestamp 1018054153
transform 1 0 4016 0 1 3280
box -16 -6 32 210
use FILL  FILL_6551
timestamp 1018054153
transform 1 0 4032 0 1 3280
box -16 -6 32 210
use FILL  FILL_6553
timestamp 1018054153
transform 1 0 4048 0 1 3280
box -16 -6 32 210
use FILL  FILL_6555
timestamp 1018054153
transform 1 0 4064 0 1 3280
box -16 -6 32 210
use FILL  FILL_6557
timestamp 1018054153
transform 1 0 4080 0 1 3280
box -16 -6 32 210
use FILL  FILL_6559
timestamp 1018054153
transform 1 0 4096 0 1 3280
box -16 -6 32 210
use FILL  FILL_6561
timestamp 1018054153
transform 1 0 4112 0 1 3280
box -16 -6 32 210
use FILL  FILL_6563
timestamp 1018054153
transform 1 0 4128 0 1 3280
box -16 -6 32 210
use FILL  FILL_6565
timestamp 1018054153
transform 1 0 4144 0 1 3280
box -16 -6 32 210
use FILL  FILL_6567
timestamp 1018054153
transform 1 0 4160 0 1 3280
box -16 -6 32 210
use FILL  FILL_6569
timestamp 1018054153
transform 1 0 4176 0 1 3280
box -16 -6 32 210
use FILL  FILL_6571
timestamp 1018054153
transform 1 0 4192 0 1 3280
box -16 -6 32 210
use FILL  FILL_6573
timestamp 1018054153
transform 1 0 4208 0 1 3280
box -16 -6 32 210
use FILL  FILL_6575
timestamp 1018054153
transform 1 0 4224 0 1 3280
box -16 -6 32 210
use FILL  FILL_6577
timestamp 1018054153
transform 1 0 4240 0 1 3280
box -16 -6 32 210
use FILL  FILL_6579
timestamp 1018054153
transform 1 0 4256 0 1 3280
box -16 -6 32 210
use FILL  FILL_6581
timestamp 1018054153
transform 1 0 4272 0 1 3280
box -16 -6 32 210
use FILL  FILL_6583
timestamp 1018054153
transform 1 0 4288 0 1 3280
box -16 -6 32 210
use FILL  FILL_6585
timestamp 1018054153
transform 1 0 4304 0 1 3280
box -16 -6 32 210
use FILL  FILL_6587
timestamp 1018054153
transform 1 0 4320 0 1 3280
box -16 -6 32 210
use FILL  FILL_6589
timestamp 1018054153
transform 1 0 4336 0 1 3280
box -16 -6 32 210
use FILL  FILL_6591
timestamp 1018054153
transform 1 0 4352 0 1 3280
box -16 -6 32 210
use FILL  FILL_6593
timestamp 1018054153
transform 1 0 4368 0 1 3280
box -16 -6 32 210
use FILL  FILL_6595
timestamp 1018054153
transform 1 0 4384 0 1 3280
box -16 -6 32 210
use FILL  FILL_6597
timestamp 1018054153
transform 1 0 4400 0 1 3280
box -16 -6 32 210
use FILL  FILL_6599
timestamp 1018054153
transform 1 0 4416 0 1 3280
box -16 -6 32 210
use FILL  FILL_6601
timestamp 1018054153
transform 1 0 4432 0 1 3280
box -16 -6 32 210
use FILL  FILL_6603
timestamp 1018054153
transform 1 0 4448 0 1 3280
box -16 -6 32 210
use FILL  FILL_6605
timestamp 1018054153
transform 1 0 4464 0 1 3280
box -16 -6 32 210
use FILL  FILL_6607
timestamp 1018054153
transform 1 0 4480 0 1 3280
box -16 -6 32 210
use FILL  FILL_6609
timestamp 1018054153
transform 1 0 4496 0 1 3280
box -16 -6 32 210
use FILL  FILL_6611
timestamp 1018054153
transform 1 0 4512 0 1 3280
box -16 -6 32 210
use FILL  FILL_6613
timestamp 1018054153
transform 1 0 4528 0 1 3280
box -16 -6 32 210
use FILL  FILL_6615
timestamp 1018054153
transform 1 0 4544 0 1 3280
box -16 -6 32 210
use FILL  FILL_6617
timestamp 1018054153
transform 1 0 4560 0 1 3280
box -16 -6 32 210
use FILL  FILL_6619
timestamp 1018054153
transform 1 0 4576 0 1 3280
box -16 -6 32 210
use FILL  FILL_6621
timestamp 1018054153
transform 1 0 4592 0 1 3280
box -16 -6 32 210
use FILL  FILL_6623
timestamp 1018054153
transform 1 0 4608 0 1 3280
box -16 -6 32 210
use FILL  FILL_6625
timestamp 1018054153
transform 1 0 4624 0 1 3280
box -16 -6 32 210
use FILL  FILL_6627
timestamp 1018054153
transform 1 0 4640 0 1 3280
box -16 -6 32 210
use FILL  FILL_6629
timestamp 1018054153
transform 1 0 4656 0 1 3280
box -16 -6 32 210
use FILL  FILL_6631
timestamp 1018054153
transform 1 0 4672 0 1 3280
box -16 -6 32 210
use FILL  FILL_6633
timestamp 1018054153
transform 1 0 4688 0 1 3280
box -16 -6 32 210
use FILL  FILL_6635
timestamp 1018054153
transform 1 0 4704 0 1 3280
box -16 -6 32 210
use FILL  FILL_6637
timestamp 1018054153
transform 1 0 4720 0 1 3280
box -16 -6 32 210
use FILL  FILL_6639
timestamp 1018054153
transform 1 0 4736 0 1 3280
box -16 -6 32 210
use FILL  FILL_6641
timestamp 1018054153
transform 1 0 4752 0 1 3280
box -16 -6 32 210
use FILL  FILL_6643
timestamp 1018054153
transform 1 0 4768 0 1 3280
box -16 -6 32 210
use FILL  FILL_6645
timestamp 1018054153
transform 1 0 4784 0 1 3280
box -16 -6 32 210
use FILL  FILL_6647
timestamp 1018054153
transform 1 0 4800 0 1 3280
box -16 -6 32 210
use FILL  FILL_6649
timestamp 1018054153
transform 1 0 4816 0 1 3280
box -16 -6 32 210
use FILL  FILL_6651
timestamp 1018054153
transform 1 0 4832 0 1 3280
box -16 -6 32 210
use FILL  FILL_6653
timestamp 1018054153
transform 1 0 4848 0 1 3280
box -16 -6 32 210
use FILL  FILL_6655
timestamp 1018054153
transform 1 0 4864 0 1 3280
box -16 -6 32 210
use FILL  FILL_6657
timestamp 1018054153
transform 1 0 4880 0 1 3280
box -16 -6 32 210
use FILL  FILL_6659
timestamp 1018054153
transform 1 0 4896 0 1 3280
box -16 -6 32 210
use FILL  FILL_6661
timestamp 1018054153
transform 1 0 4912 0 1 3280
box -16 -6 32 210
use FILL  FILL_6663
timestamp 1018054153
transform 1 0 4928 0 1 3280
box -16 -6 32 210
use FILL  FILL_6665
timestamp 1018054153
transform 1 0 4944 0 1 3280
box -16 -6 32 210
use FILL  FILL_6667
timestamp 1018054153
transform 1 0 4960 0 1 3280
box -16 -6 32 210
use FILL  FILL_6669
timestamp 1018054153
transform 1 0 4976 0 1 3280
box -16 -6 32 210
use FILL  FILL_6671
timestamp 1018054153
transform 1 0 4992 0 1 3280
box -16 -6 32 210
use FILL  FILL_6673
timestamp 1018054153
transform 1 0 5008 0 1 3280
box -16 -6 32 210
use FILL  FILL_6675
timestamp 1018054153
transform 1 0 5024 0 1 3280
box -16 -6 32 210
use FILL  FILL_6677
timestamp 1018054153
transform 1 0 5040 0 1 3280
box -16 -6 32 210
use FILL  FILL_6679
timestamp 1018054153
transform 1 0 5056 0 1 3280
box -16 -6 32 210
use FILL  FILL_6681
timestamp 1018054153
transform 1 0 5072 0 1 3280
box -16 -6 32 210
use FILL  FILL_6683
timestamp 1018054153
transform 1 0 5088 0 1 3280
box -16 -6 32 210
use FILL  FILL_6685
timestamp 1018054153
transform 1 0 5104 0 1 3280
box -16 -6 32 210
use FILL  FILL_6687
timestamp 1018054153
transform 1 0 5120 0 1 3280
box -16 -6 32 210
use FILL  FILL_6689
timestamp 1018054153
transform 1 0 5136 0 1 3280
box -16 -6 32 210
use FILL  FILL_6691
timestamp 1018054153
transform 1 0 5152 0 1 3280
box -16 -6 32 210
use FILL  FILL_6693
timestamp 1018054153
transform 1 0 5168 0 1 3280
box -16 -6 32 210
use FILL  FILL_6695
timestamp 1018054153
transform 1 0 5184 0 1 3280
box -16 -6 32 210
use FILL  FILL_6697
timestamp 1018054153
transform 1 0 5200 0 1 3280
box -16 -6 32 210
use FILL  FILL_6699
timestamp 1018054153
transform 1 0 5216 0 1 3280
box -16 -6 32 210
use FILL  FILL_6701
timestamp 1018054153
transform 1 0 5232 0 1 3280
box -16 -6 32 210
use FILL  FILL_6703
timestamp 1018054153
transform 1 0 5248 0 1 3280
box -16 -6 32 210
use FILL  FILL_6705
timestamp 1018054153
transform 1 0 5264 0 1 3280
box -16 -6 32 210
use FILL  FILL_6707
timestamp 1018054153
transform 1 0 5280 0 1 3280
box -16 -6 32 210
use FILL  FILL_6709
timestamp 1018054153
transform 1 0 5296 0 1 3280
box -16 -6 32 210
use FILL  FILL_6711
timestamp 1018054153
transform 1 0 5312 0 1 3280
box -16 -6 32 210
use FILL  FILL_6713
timestamp 1018054153
transform 1 0 5328 0 1 3280
box -16 -6 32 210
use FILL  FILL_6715
timestamp 1018054153
transform 1 0 5344 0 1 3280
box -16 -6 32 210
use FILL  FILL_6717
timestamp 1018054153
transform 1 0 5360 0 1 3280
box -16 -6 32 210
use FILL  FILL_6719
timestamp 1018054153
transform 1 0 5376 0 1 3280
box -16 -6 32 210
use FILL  FILL_6721
timestamp 1018054153
transform 1 0 5392 0 1 3280
box -16 -6 32 210
use FILL  FILL_6723
timestamp 1018054153
transform 1 0 5408 0 1 3280
box -16 -6 32 210
use FILL  FILL_6725
timestamp 1018054153
transform 1 0 5424 0 1 3280
box -16 -6 32 210
use FILL  FILL_6727
timestamp 1018054153
transform 1 0 5440 0 1 3280
box -16 -6 32 210
use FILL  FILL_6729
timestamp 1018054153
transform 1 0 5456 0 1 3280
box -16 -6 32 210
use FILL  FILL_6731
timestamp 1018054153
transform 1 0 5472 0 1 3280
box -16 -6 32 210
use FILL  FILL_6733
timestamp 1018054153
transform 1 0 5488 0 1 3280
box -16 -6 32 210
use FILL  FILL_6735
timestamp 1018054153
transform 1 0 5504 0 1 3280
box -16 -6 32 210
use FILL  FILL_6737
timestamp 1018054153
transform 1 0 5520 0 1 3280
box -16 -6 32 210
use FILL  FILL_6739
timestamp 1018054153
transform 1 0 5536 0 1 3280
box -16 -6 32 210
use FILL  FILL_6741
timestamp 1018054153
transform 1 0 5552 0 1 3280
box -16 -6 32 210
use FILL  FILL_6743
timestamp 1018054153
transform 1 0 5568 0 1 3280
box -16 -6 32 210
use FILL  FILL_6745
timestamp 1018054153
transform 1 0 5584 0 1 3280
box -16 -6 32 210
use FILL  FILL_6747
timestamp 1018054153
transform 1 0 5600 0 1 3280
box -16 -6 32 210
use FILL  FILL_6749
timestamp 1018054153
transform 1 0 5616 0 1 3280
box -16 -6 32 210
use FILL  FILL_6751
timestamp 1018054153
transform 1 0 5632 0 1 3280
box -16 -6 32 210
use FILL  FILL_6753
timestamp 1018054153
transform 1 0 5648 0 1 3280
box -16 -6 32 210
use FILL  FILL_6755
timestamp 1018054153
transform 1 0 5664 0 1 3280
box -16 -6 32 210
use FILL  FILL_6757
timestamp 1018054153
transform 1 0 5680 0 1 3280
box -16 -6 32 210
use FILL  FILL_6759
timestamp 1018054153
transform 1 0 5696 0 1 3280
box -16 -6 32 210
use FILL  FILL_6761
timestamp 1018054153
transform 1 0 5712 0 1 3280
box -16 -6 32 210
use FILL  FILL_6763
timestamp 1018054153
transform 1 0 5728 0 1 3280
box -16 -6 32 210
use FILL  FILL_6765
timestamp 1018054153
transform 1 0 5744 0 1 3280
box -16 -6 32 210
use FILL  FILL_6767
timestamp 1018054153
transform 1 0 5760 0 1 3280
box -16 -6 32 210
use FILL  FILL_6769
timestamp 1018054153
transform 1 0 5776 0 1 3280
box -16 -6 32 210
use FILL  FILL_6771
timestamp 1018054153
transform 1 0 5792 0 1 3280
box -16 -6 32 210
use FILL  FILL_6773
timestamp 1018054153
transform 1 0 5808 0 1 3280
box -16 -6 32 210
use FILL  FILL_6775
timestamp 1018054153
transform 1 0 5824 0 1 3280
box -16 -6 32 210
use FILL  FILL_6777
timestamp 1018054153
transform 1 0 5840 0 1 3280
box -16 -6 32 210
use FILL  FILL_6779
timestamp 1018054153
transform 1 0 5856 0 1 3280
box -16 -6 32 210
use FILL  FILL_6781
timestamp 1018054153
transform 1 0 5872 0 1 3280
box -16 -6 32 210
use FILL  FILL_6783
timestamp 1018054153
transform 1 0 5888 0 1 3280
box -16 -6 32 210
use FILL  FILL_6785
timestamp 1018054153
transform 1 0 5904 0 1 3280
box -16 -6 32 210
use FILL  FILL_6787
timestamp 1018054153
transform 1 0 5920 0 1 3280
box -16 -6 32 210
use FILL  FILL_6789
timestamp 1018054153
transform 1 0 5936 0 1 3280
box -16 -6 32 210
use FILL  FILL_6791
timestamp 1018054153
transform 1 0 5952 0 1 3280
box -16 -6 32 210
use FILL  FILL_6793
timestamp 1018054153
transform 1 0 5968 0 1 3280
box -16 -6 32 210
use FILL  FILL_6795
timestamp 1018054153
transform 1 0 5984 0 1 3280
box -16 -6 32 210
use FILL  FILL_6797
timestamp 1018054153
transform 1 0 6000 0 1 3280
box -16 -6 32 210
use FILL  FILL_6799
timestamp 1018054153
transform 1 0 6016 0 1 3280
box -16 -6 32 210
use FILL  FILL_6801
timestamp 1018054153
transform 1 0 6032 0 1 3280
box -16 -6 32 210
use FILL  FILL_6803
timestamp 1018054153
transform 1 0 6048 0 1 3280
box -16 -6 32 210
use FILL  FILL_6805
timestamp 1018054153
transform 1 0 6064 0 1 3280
box -16 -6 32 210
use FILL  FILL_6807
timestamp 1018054153
transform 1 0 6080 0 1 3280
box -16 -6 32 210
use FILL  FILL_6809
timestamp 1018054153
transform 1 0 6096 0 1 3280
box -16 -6 32 210
use FILL  FILL_6811
timestamp 1018054153
transform 1 0 6112 0 1 3280
box -16 -6 32 210
use FILL  FILL_6813
timestamp 1018054153
transform 1 0 6128 0 1 3280
box -16 -6 32 210
use FILL  FILL_6815
timestamp 1018054153
transform 1 0 6144 0 1 3280
box -16 -6 32 210
use FILL  FILL_6817
timestamp 1018054153
transform 1 0 6160 0 1 3280
box -16 -6 32 210
use FILL  FILL_6819
timestamp 1018054153
transform 1 0 6176 0 1 3280
box -16 -6 32 210
use FILL  FILL_6821
timestamp 1018054153
transform 1 0 6192 0 1 3280
box -16 -6 32 210
use FILL  FILL_6823
timestamp 1018054153
transform 1 0 6208 0 1 3280
box -16 -6 32 210
use FILL  FILL_6825
timestamp 1018054153
transform 1 0 6224 0 1 3280
box -16 -6 32 210
use FILL  FILL_6827
timestamp 1018054153
transform 1 0 6240 0 1 3280
box -16 -6 32 210
use FILL  FILL_6829
timestamp 1018054153
transform 1 0 6256 0 1 3280
box -16 -6 32 210
use FILL  FILL_6831
timestamp 1018054153
transform 1 0 6272 0 1 3280
box -16 -6 32 210
use FILL  FILL_6833
timestamp 1018054153
transform 1 0 6288 0 1 3280
box -16 -6 32 210
use FILL  FILL_6835
timestamp 1018054153
transform 1 0 6304 0 1 3280
box -16 -6 32 210
use FILL  FILL_6837
timestamp 1018054153
transform 1 0 6320 0 1 3280
box -16 -6 32 210
use FILL  FILL_6839
timestamp 1018054153
transform 1 0 6336 0 1 3280
box -16 -6 32 210
use FILL  FILL_6841
timestamp 1018054153
transform 1 0 6352 0 1 3280
box -16 -6 32 210
use FILL  FILL_6843
timestamp 1018054153
transform 1 0 6368 0 1 3280
box -16 -6 32 210
use FILL  FILL_6845
timestamp 1018054153
transform 1 0 6384 0 1 3280
box -16 -6 32 210
use FILL  FILL_6847
timestamp 1018054153
transform 1 0 6400 0 1 3280
box -16 -6 32 210
use FILL  FILL_6849
timestamp 1018054153
transform 1 0 6416 0 1 3280
box -16 -6 32 210
use FILL  FILL_6851
timestamp 1018054153
transform 1 0 6432 0 1 3280
box -16 -6 32 210
use FILL  FILL_6853
timestamp 1018054153
transform 1 0 6448 0 1 3280
box -16 -6 32 210
use FILL  FILL_6855
timestamp 1018054153
transform 1 0 6464 0 1 3280
box -16 -6 32 210
use FILL  FILL_6857
timestamp 1018054153
transform 1 0 6480 0 1 3280
box -16 -6 32 210
use FILL  FILL_6859
timestamp 1018054153
transform 1 0 6496 0 1 3280
box -16 -6 32 210
use FILL  FILL_6861
timestamp 1018054153
transform 1 0 6512 0 1 3280
box -16 -6 32 210
use FILL  FILL_6863
timestamp 1018054153
transform 1 0 6528 0 1 3280
box -16 -6 32 210
use FILL  FILL_6865
timestamp 1018054153
transform 1 0 6544 0 1 3280
box -16 -6 32 210
use FILL  FILL_6867
timestamp 1018054153
transform 1 0 6560 0 1 3280
box -16 -6 32 210
use FILL  FILL_6869
timestamp 1018054153
transform 1 0 6576 0 1 3280
box -16 -6 32 210
use FILL  FILL_6871
timestamp 1018054153
transform 1 0 6592 0 1 3280
box -16 -6 32 210
use FILL  FILL_6873
timestamp 1018054153
transform 1 0 6608 0 1 3280
box -16 -6 32 210
use FILL  FILL_6875
timestamp 1018054153
transform 1 0 6624 0 1 3280
box -16 -6 32 210
use FILL  FILL_6877
timestamp 1018054153
transform 1 0 6640 0 1 3280
box -16 -6 32 210
use FILL  FILL_6879
timestamp 1018054153
transform 1 0 6656 0 1 3280
box -16 -6 32 210
use FILL  FILL_6881
timestamp 1018054153
transform 1 0 6672 0 1 3280
box -16 -6 32 210
use FILL  FILL_6883
timestamp 1018054153
transform 1 0 6688 0 1 3280
box -16 -6 32 210
use FILL  FILL_6885
timestamp 1018054153
transform 1 0 6704 0 1 3280
box -16 -6 32 210
use FILL  FILL_6887
timestamp 1018054153
transform 1 0 6720 0 1 3280
box -16 -6 32 210
use FILL  FILL_6889
timestamp 1018054153
transform 1 0 6736 0 1 3280
box -16 -6 32 210
use FILL  FILL_6891
timestamp 1018054153
transform 1 0 6752 0 1 3280
box -16 -6 32 210
use FILL  FILL_6893
timestamp 1018054153
transform 1 0 6768 0 1 3280
box -16 -6 32 210
use FILL  FILL_6895
timestamp 1018054153
transform 1 0 6784 0 1 3280
box -16 -6 32 210
use FILL  FILL_6897
timestamp 1018054153
transform 1 0 6800 0 1 3280
box -16 -6 32 210
use FILL  FILL_6899
timestamp 1018054153
transform 1 0 6816 0 1 3280
box -16 -6 32 210
use FILL  FILL_6901
timestamp 1018054153
transform 1 0 6832 0 1 3280
box -16 -6 32 210
use FILL  FILL_6903
timestamp 1018054153
transform 1 0 6848 0 1 3280
box -16 -6 32 210
use FILL  FILL_6905
timestamp 1018054153
transform 1 0 6864 0 1 3280
box -16 -6 32 210
use FILL  FILL_6907
timestamp 1018054153
transform 1 0 6880 0 1 3280
box -16 -6 32 210
use FILL  FILL_6909
timestamp 1018054153
transform 1 0 6896 0 1 3280
box -16 -6 32 210
use FILL  FILL_6911
timestamp 1018054153
transform 1 0 6912 0 1 3280
box -16 -6 32 210
use FILL  FILL_6913
timestamp 1018054153
transform 1 0 6928 0 1 3280
box -16 -6 32 210
use FILL  FILL_6915
timestamp 1018054153
transform 1 0 6944 0 1 3280
box -16 -6 32 210
use FILL  FILL_6917
timestamp 1018054153
transform 1 0 6960 0 1 3280
box -16 -6 32 210
use FILL  FILL_6919
timestamp 1018054153
transform 1 0 6976 0 1 3280
box -16 -6 32 210
use FILL  FILL_6921
timestamp 1018054153
transform 1 0 6992 0 1 3280
box -16 -6 32 210
use FILL  FILL_6923
timestamp 1018054153
transform 1 0 7008 0 1 3280
box -16 -6 32 210
use FILL  FILL_6925
timestamp 1018054153
transform 1 0 7024 0 1 3280
box -16 -6 32 210
use FILL  FILL_6927
timestamp 1018054153
transform 1 0 7040 0 1 3280
box -16 -6 32 210
use FILL  FILL_6929
timestamp 1018054153
transform 1 0 7056 0 1 3280
box -16 -6 32 210
use FILL  FILL_6931
timestamp 1018054153
transform 1 0 7072 0 1 3280
box -16 -6 32 210
use FILL  FILL_6933
timestamp 1018054153
transform 1 0 7088 0 1 3280
box -16 -6 32 210
use FILL  FILL_6935
timestamp 1018054153
transform 1 0 7104 0 1 3280
box -16 -6 32 210
use FILL  FILL_6937
timestamp 1018054153
transform 1 0 7120 0 1 3280
box -16 -6 32 210
use FILL  FILL_6939
timestamp 1018054153
transform 1 0 7136 0 1 3280
box -16 -6 32 210
use FILL  FILL_6941
timestamp 1018054153
transform 1 0 7152 0 1 3280
box -16 -6 32 210
use FILL  FILL_6943
timestamp 1018054153
transform 1 0 7168 0 1 3280
box -16 -6 32 210
use FILL  FILL_6945
timestamp 1018054153
transform 1 0 7184 0 1 3280
box -16 -6 32 210
use FILL  FILL_6947
timestamp 1018054153
transform 1 0 7200 0 1 3280
box -16 -6 32 210
use FILL  FILL_6949
timestamp 1018054153
transform 1 0 7216 0 1 3280
box -16 -6 32 210
use FILL  FILL_6951
timestamp 1018054153
transform 1 0 7232 0 1 3280
box -16 -6 32 210
use FILL  FILL_6953
timestamp 1018054153
transform 1 0 7248 0 1 3280
box -16 -6 32 210
use FILL  FILL_6955
timestamp 1018054153
transform 1 0 7264 0 1 3280
box -16 -6 32 210
use FILL  FILL_6957
timestamp 1018054153
transform 1 0 7280 0 1 3280
box -16 -6 32 210
use FILL  FILL_6959
timestamp 1018054153
transform 1 0 7296 0 1 3280
box -16 -6 32 210
use FILL  FILL_6961
timestamp 1018054153
transform 1 0 7312 0 1 3280
box -16 -6 32 210
use FILL  FILL_6963
timestamp 1018054153
transform 1 0 7328 0 1 3280
box -16 -6 32 210
use FILL  FILL_6965
timestamp 1018054153
transform 1 0 7344 0 1 3280
box -16 -6 32 210
use FILL  FILL_6967
timestamp 1018054153
transform 1 0 7360 0 1 3280
box -16 -6 32 210
use FILL  FILL_6969
timestamp 1018054153
transform 1 0 7376 0 1 3280
box -16 -6 32 210
use FILL  FILL_6971
timestamp 1018054153
transform 1 0 7392 0 1 3280
box -16 -6 32 210
use FILL  FILL_6973
timestamp 1018054153
transform 1 0 7408 0 1 3280
box -16 -6 32 210
use FILL  FILL_6975
timestamp 1018054153
transform 1 0 7424 0 1 3280
box -16 -6 32 210
use FILL  FILL_6977
timestamp 1018054153
transform 1 0 7440 0 1 3280
box -16 -6 32 210
use FILL  FILL_6979
timestamp 1018054153
transform 1 0 7456 0 1 3280
box -16 -6 32 210
use FILL  FILL_6981
timestamp 1018054153
transform 1 0 7472 0 1 3280
box -16 -6 32 210
use FILL  FILL_6983
timestamp 1018054153
transform 1 0 7488 0 1 3280
box -16 -6 32 210
use FILL  FILL_6985
timestamp 1018054153
transform 1 0 7504 0 1 3280
box -16 -6 32 210
use FILL  FILL_6987
timestamp 1018054153
transform 1 0 7520 0 1 3280
box -16 -6 32 210
use FILL  FILL_6989
timestamp 1018054153
transform 1 0 7536 0 1 3280
box -16 -6 32 210
use FILL  FILL_6991
timestamp 1018054153
transform 1 0 7552 0 1 3280
box -16 -6 32 210
use FILL  FILL_6993
timestamp 1018054153
transform 1 0 7568 0 1 3280
box -16 -6 32 210
use FILL  FILL_6995
timestamp 1018054153
transform 1 0 7584 0 1 3280
box -16 -6 32 210
use FILL  FILL_6997
timestamp 1018054153
transform 1 0 7600 0 1 3280
box -16 -6 32 210
use FILL  FILL_6999
timestamp 1018054153
transform 1 0 7616 0 1 3280
box -16 -6 32 210
use FILL  FILL_7001
timestamp 1018054153
transform 1 0 7632 0 1 3280
box -16 -6 32 210
use FILL  FILL_7003
timestamp 1018054153
transform 1 0 7648 0 1 3280
box -16 -6 32 210
use FILL  FILL_7005
timestamp 1018054153
transform 1 0 7664 0 1 3280
box -16 -6 32 210
use FILL  FILL_7007
timestamp 1018054153
transform 1 0 7680 0 1 3280
box -16 -6 32 210
use FILL  FILL_7009
timestamp 1018054153
transform 1 0 7696 0 1 3280
box -16 -6 32 210
use FILL  FILL_7011
timestamp 1018054153
transform 1 0 7712 0 1 3280
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_41
timestamp 1542725905
transform 1 0 7908 0 1 3280
box -48 -6 48 6
use PADINC  PADINC_9
timestamp 1084294328
transform 0 -1 2000 1 0 3200
box -12 -6 606 2000
use M2_M1  M2_M1_286
timestamp 1542725905
transform 1 0 6296 0 1 3170
box -4 -4 4 4
use PADOUT  PADOUT_3
timestamp 1084294529
transform 0 1 8000 -1 0 3800
box -12 -6 606 2000
use M2_M1  M2_M1_287
timestamp 1542725905
transform 1 0 7976 0 1 3170
box -4 -4 4 4
use M3_M2  M3_M2_124
timestamp 1542725905
transform 1 0 7976 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_125
timestamp 1542725905
transform 1 0 8002 0 1 3110
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_42
timestamp 1542725905
transform 1 0 2212 0 1 3080
box -48 -6 48 6
use FILL  FILL_6332
timestamp 1018054153
transform 1 0 2272 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6334
timestamp 1018054153
transform 1 0 2288 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6336
timestamp 1018054153
transform 1 0 2304 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6338
timestamp 1018054153
transform 1 0 2320 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6340
timestamp 1018054153
transform 1 0 2336 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6342
timestamp 1018054153
transform 1 0 2352 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6344
timestamp 1018054153
transform 1 0 2368 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6346
timestamp 1018054153
transform 1 0 2384 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6348
timestamp 1018054153
transform 1 0 2400 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6350
timestamp 1018054153
transform 1 0 2416 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6352
timestamp 1018054153
transform 1 0 2432 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6354
timestamp 1018054153
transform 1 0 2448 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6356
timestamp 1018054153
transform 1 0 2464 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6358
timestamp 1018054153
transform 1 0 2480 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6360
timestamp 1018054153
transform 1 0 2496 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6362
timestamp 1018054153
transform 1 0 2512 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6364
timestamp 1018054153
transform 1 0 2528 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6366
timestamp 1018054153
transform 1 0 2544 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6368
timestamp 1018054153
transform 1 0 2560 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6370
timestamp 1018054153
transform 1 0 2576 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6372
timestamp 1018054153
transform 1 0 2592 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6374
timestamp 1018054153
transform 1 0 2608 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6376
timestamp 1018054153
transform 1 0 2624 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6378
timestamp 1018054153
transform 1 0 2640 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6380
timestamp 1018054153
transform 1 0 2656 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6382
timestamp 1018054153
transform 1 0 2672 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6384
timestamp 1018054153
transform 1 0 2688 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6386
timestamp 1018054153
transform 1 0 2704 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6388
timestamp 1018054153
transform 1 0 2720 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6390
timestamp 1018054153
transform 1 0 2736 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6392
timestamp 1018054153
transform 1 0 2752 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6394
timestamp 1018054153
transform 1 0 2768 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6396
timestamp 1018054153
transform 1 0 2784 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6398
timestamp 1018054153
transform 1 0 2800 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6400
timestamp 1018054153
transform 1 0 2816 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6402
timestamp 1018054153
transform 1 0 2832 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6404
timestamp 1018054153
transform 1 0 2848 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6406
timestamp 1018054153
transform 1 0 2864 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6408
timestamp 1018054153
transform 1 0 2880 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6410
timestamp 1018054153
transform 1 0 2896 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6412
timestamp 1018054153
transform 1 0 2912 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6414
timestamp 1018054153
transform 1 0 2928 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6416
timestamp 1018054153
transform 1 0 2944 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6418
timestamp 1018054153
transform 1 0 2960 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6420
timestamp 1018054153
transform 1 0 2976 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6422
timestamp 1018054153
transform 1 0 2992 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6424
timestamp 1018054153
transform 1 0 3008 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6426
timestamp 1018054153
transform 1 0 3024 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6428
timestamp 1018054153
transform 1 0 3040 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6430
timestamp 1018054153
transform 1 0 3056 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6432
timestamp 1018054153
transform 1 0 3072 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6434
timestamp 1018054153
transform 1 0 3088 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6436
timestamp 1018054153
transform 1 0 3104 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6438
timestamp 1018054153
transform 1 0 3120 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6440
timestamp 1018054153
transform 1 0 3136 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6442
timestamp 1018054153
transform 1 0 3152 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6444
timestamp 1018054153
transform 1 0 3168 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6446
timestamp 1018054153
transform 1 0 3184 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6448
timestamp 1018054153
transform 1 0 3200 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6450
timestamp 1018054153
transform 1 0 3216 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6452
timestamp 1018054153
transform 1 0 3232 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6454
timestamp 1018054153
transform 1 0 3248 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6456
timestamp 1018054153
transform 1 0 3264 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6458
timestamp 1018054153
transform 1 0 3280 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6460
timestamp 1018054153
transform 1 0 3296 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6462
timestamp 1018054153
transform 1 0 3312 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6464
timestamp 1018054153
transform 1 0 3328 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6466
timestamp 1018054153
transform 1 0 3344 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6468
timestamp 1018054153
transform 1 0 3360 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6470
timestamp 1018054153
transform 1 0 3376 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6472
timestamp 1018054153
transform 1 0 3392 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6474
timestamp 1018054153
transform 1 0 3408 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6476
timestamp 1018054153
transform 1 0 3424 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6478
timestamp 1018054153
transform 1 0 3440 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6480
timestamp 1018054153
transform 1 0 3456 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6482
timestamp 1018054153
transform 1 0 3472 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6484
timestamp 1018054153
transform 1 0 3488 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6486
timestamp 1018054153
transform 1 0 3504 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6488
timestamp 1018054153
transform 1 0 3520 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6490
timestamp 1018054153
transform 1 0 3536 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6492
timestamp 1018054153
transform 1 0 3552 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6494
timestamp 1018054153
transform 1 0 3568 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6496
timestamp 1018054153
transform 1 0 3584 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6498
timestamp 1018054153
transform 1 0 3600 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6500
timestamp 1018054153
transform 1 0 3616 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6502
timestamp 1018054153
transform 1 0 3632 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6504
timestamp 1018054153
transform 1 0 3648 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6506
timestamp 1018054153
transform 1 0 3664 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6508
timestamp 1018054153
transform 1 0 3680 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6510
timestamp 1018054153
transform 1 0 3696 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6512
timestamp 1018054153
transform 1 0 3712 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6514
timestamp 1018054153
transform 1 0 3728 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6516
timestamp 1018054153
transform 1 0 3744 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6518
timestamp 1018054153
transform 1 0 3760 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6520
timestamp 1018054153
transform 1 0 3776 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6522
timestamp 1018054153
transform 1 0 3792 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6524
timestamp 1018054153
transform 1 0 3808 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6526
timestamp 1018054153
transform 1 0 3824 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6528
timestamp 1018054153
transform 1 0 3840 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6530
timestamp 1018054153
transform 1 0 3856 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6532
timestamp 1018054153
transform 1 0 3872 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6534
timestamp 1018054153
transform 1 0 3888 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6536
timestamp 1018054153
transform 1 0 3904 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6538
timestamp 1018054153
transform 1 0 3920 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6540
timestamp 1018054153
transform 1 0 3936 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6542
timestamp 1018054153
transform 1 0 3952 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6544
timestamp 1018054153
transform 1 0 3968 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6546
timestamp 1018054153
transform 1 0 3984 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6548
timestamp 1018054153
transform 1 0 4000 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6550
timestamp 1018054153
transform 1 0 4016 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6552
timestamp 1018054153
transform 1 0 4032 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6554
timestamp 1018054153
transform 1 0 4048 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6556
timestamp 1018054153
transform 1 0 4064 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6558
timestamp 1018054153
transform 1 0 4080 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6560
timestamp 1018054153
transform 1 0 4096 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6562
timestamp 1018054153
transform 1 0 4112 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6564
timestamp 1018054153
transform 1 0 4128 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6566
timestamp 1018054153
transform 1 0 4144 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6568
timestamp 1018054153
transform 1 0 4160 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6570
timestamp 1018054153
transform 1 0 4176 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6572
timestamp 1018054153
transform 1 0 4192 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6574
timestamp 1018054153
transform 1 0 4208 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6576
timestamp 1018054153
transform 1 0 4224 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6578
timestamp 1018054153
transform 1 0 4240 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6580
timestamp 1018054153
transform 1 0 4256 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6582
timestamp 1018054153
transform 1 0 4272 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6584
timestamp 1018054153
transform 1 0 4288 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6586
timestamp 1018054153
transform 1 0 4304 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6588
timestamp 1018054153
transform 1 0 4320 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6590
timestamp 1018054153
transform 1 0 4336 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6592
timestamp 1018054153
transform 1 0 4352 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6594
timestamp 1018054153
transform 1 0 4368 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6596
timestamp 1018054153
transform 1 0 4384 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6598
timestamp 1018054153
transform 1 0 4400 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6600
timestamp 1018054153
transform 1 0 4416 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6602
timestamp 1018054153
transform 1 0 4432 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6604
timestamp 1018054153
transform 1 0 4448 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6606
timestamp 1018054153
transform 1 0 4464 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6608
timestamp 1018054153
transform 1 0 4480 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6610
timestamp 1018054153
transform 1 0 4496 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6612
timestamp 1018054153
transform 1 0 4512 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6614
timestamp 1018054153
transform 1 0 4528 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6616
timestamp 1018054153
transform 1 0 4544 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6618
timestamp 1018054153
transform 1 0 4560 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6620
timestamp 1018054153
transform 1 0 4576 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6622
timestamp 1018054153
transform 1 0 4592 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6624
timestamp 1018054153
transform 1 0 4608 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6626
timestamp 1018054153
transform 1 0 4624 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6628
timestamp 1018054153
transform 1 0 4640 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6630
timestamp 1018054153
transform 1 0 4656 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6632
timestamp 1018054153
transform 1 0 4672 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6634
timestamp 1018054153
transform 1 0 4688 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6636
timestamp 1018054153
transform 1 0 4704 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6638
timestamp 1018054153
transform 1 0 4720 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6640
timestamp 1018054153
transform 1 0 4736 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6642
timestamp 1018054153
transform 1 0 4752 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6644
timestamp 1018054153
transform 1 0 4768 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6646
timestamp 1018054153
transform 1 0 4784 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6648
timestamp 1018054153
transform 1 0 4800 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6650
timestamp 1018054153
transform 1 0 4816 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6652
timestamp 1018054153
transform 1 0 4832 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6654
timestamp 1018054153
transform 1 0 4848 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6656
timestamp 1018054153
transform 1 0 4864 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6658
timestamp 1018054153
transform 1 0 4880 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6660
timestamp 1018054153
transform 1 0 4896 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6662
timestamp 1018054153
transform 1 0 4912 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6664
timestamp 1018054153
transform 1 0 4928 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6666
timestamp 1018054153
transform 1 0 4944 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6668
timestamp 1018054153
transform 1 0 4960 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6670
timestamp 1018054153
transform 1 0 4976 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6672
timestamp 1018054153
transform 1 0 4992 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6674
timestamp 1018054153
transform 1 0 5008 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6676
timestamp 1018054153
transform 1 0 5024 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6678
timestamp 1018054153
transform 1 0 5040 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6680
timestamp 1018054153
transform 1 0 5056 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6682
timestamp 1018054153
transform 1 0 5072 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6684
timestamp 1018054153
transform 1 0 5088 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6686
timestamp 1018054153
transform 1 0 5104 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6688
timestamp 1018054153
transform 1 0 5120 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6690
timestamp 1018054153
transform 1 0 5136 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6692
timestamp 1018054153
transform 1 0 5152 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6694
timestamp 1018054153
transform 1 0 5168 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6696
timestamp 1018054153
transform 1 0 5184 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6698
timestamp 1018054153
transform 1 0 5200 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6700
timestamp 1018054153
transform 1 0 5216 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6702
timestamp 1018054153
transform 1 0 5232 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6704
timestamp 1018054153
transform 1 0 5248 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6706
timestamp 1018054153
transform 1 0 5264 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6708
timestamp 1018054153
transform 1 0 5280 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6710
timestamp 1018054153
transform 1 0 5296 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6712
timestamp 1018054153
transform 1 0 5312 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6714
timestamp 1018054153
transform 1 0 5328 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6716
timestamp 1018054153
transform 1 0 5344 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6718
timestamp 1018054153
transform 1 0 5360 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6720
timestamp 1018054153
transform 1 0 5376 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6722
timestamp 1018054153
transform 1 0 5392 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6724
timestamp 1018054153
transform 1 0 5408 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6726
timestamp 1018054153
transform 1 0 5424 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6728
timestamp 1018054153
transform 1 0 5440 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6730
timestamp 1018054153
transform 1 0 5456 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6732
timestamp 1018054153
transform 1 0 5472 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6734
timestamp 1018054153
transform 1 0 5488 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6736
timestamp 1018054153
transform 1 0 5504 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6738
timestamp 1018054153
transform 1 0 5520 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6740
timestamp 1018054153
transform 1 0 5536 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6742
timestamp 1018054153
transform 1 0 5552 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6744
timestamp 1018054153
transform 1 0 5568 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6746
timestamp 1018054153
transform 1 0 5584 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6748
timestamp 1018054153
transform 1 0 5600 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6750
timestamp 1018054153
transform 1 0 5616 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6752
timestamp 1018054153
transform 1 0 5632 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6754
timestamp 1018054153
transform 1 0 5648 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6756
timestamp 1018054153
transform 1 0 5664 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6758
timestamp 1018054153
transform 1 0 5680 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6760
timestamp 1018054153
transform 1 0 5696 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6762
timestamp 1018054153
transform 1 0 5712 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6764
timestamp 1018054153
transform 1 0 5728 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6766
timestamp 1018054153
transform 1 0 5744 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6768
timestamp 1018054153
transform 1 0 5760 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6770
timestamp 1018054153
transform 1 0 5776 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6772
timestamp 1018054153
transform 1 0 5792 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6774
timestamp 1018054153
transform 1 0 5808 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6776
timestamp 1018054153
transform 1 0 5824 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6778
timestamp 1018054153
transform 1 0 5840 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6780
timestamp 1018054153
transform 1 0 5856 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6782
timestamp 1018054153
transform 1 0 5872 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6784
timestamp 1018054153
transform 1 0 5888 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6786
timestamp 1018054153
transform 1 0 5904 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6788
timestamp 1018054153
transform 1 0 5920 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6790
timestamp 1018054153
transform 1 0 5936 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6792
timestamp 1018054153
transform 1 0 5952 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6794
timestamp 1018054153
transform 1 0 5968 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6796
timestamp 1018054153
transform 1 0 5984 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6798
timestamp 1018054153
transform 1 0 6000 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6800
timestamp 1018054153
transform 1 0 6016 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6802
timestamp 1018054153
transform 1 0 6032 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6804
timestamp 1018054153
transform 1 0 6048 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6806
timestamp 1018054153
transform 1 0 6064 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6808
timestamp 1018054153
transform 1 0 6080 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6810
timestamp 1018054153
transform 1 0 6096 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6812
timestamp 1018054153
transform 1 0 6112 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6814
timestamp 1018054153
transform 1 0 6128 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6816
timestamp 1018054153
transform 1 0 6144 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6818
timestamp 1018054153
transform 1 0 6160 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6820
timestamp 1018054153
transform 1 0 6176 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6822
timestamp 1018054153
transform 1 0 6192 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6824
timestamp 1018054153
transform 1 0 6208 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6826
timestamp 1018054153
transform 1 0 6224 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6828
timestamp 1018054153
transform 1 0 6240 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6830
timestamp 1018054153
transform 1 0 6256 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6832
timestamp 1018054153
transform 1 0 6272 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6834
timestamp 1018054153
transform 1 0 6288 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6836
timestamp 1018054153
transform 1 0 6304 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6838
timestamp 1018054153
transform 1 0 6320 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6840
timestamp 1018054153
transform 1 0 6336 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6842
timestamp 1018054153
transform 1 0 6352 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6844
timestamp 1018054153
transform 1 0 6368 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6846
timestamp 1018054153
transform 1 0 6384 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6848
timestamp 1018054153
transform 1 0 6400 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6850
timestamp 1018054153
transform 1 0 6416 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6852
timestamp 1018054153
transform 1 0 6432 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6854
timestamp 1018054153
transform 1 0 6448 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6856
timestamp 1018054153
transform 1 0 6464 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6858
timestamp 1018054153
transform 1 0 6480 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6860
timestamp 1018054153
transform 1 0 6496 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6862
timestamp 1018054153
transform 1 0 6512 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6864
timestamp 1018054153
transform 1 0 6528 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6866
timestamp 1018054153
transform 1 0 6544 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6868
timestamp 1018054153
transform 1 0 6560 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6870
timestamp 1018054153
transform 1 0 6576 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6872
timestamp 1018054153
transform 1 0 6592 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6874
timestamp 1018054153
transform 1 0 6608 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6876
timestamp 1018054153
transform 1 0 6624 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6878
timestamp 1018054153
transform 1 0 6640 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6880
timestamp 1018054153
transform 1 0 6656 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6882
timestamp 1018054153
transform 1 0 6672 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6884
timestamp 1018054153
transform 1 0 6688 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6886
timestamp 1018054153
transform 1 0 6704 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6888
timestamp 1018054153
transform 1 0 6720 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6890
timestamp 1018054153
transform 1 0 6736 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6892
timestamp 1018054153
transform 1 0 6752 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6894
timestamp 1018054153
transform 1 0 6768 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6896
timestamp 1018054153
transform 1 0 6784 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6898
timestamp 1018054153
transform 1 0 6800 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6900
timestamp 1018054153
transform 1 0 6816 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6902
timestamp 1018054153
transform 1 0 6832 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6904
timestamp 1018054153
transform 1 0 6848 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6906
timestamp 1018054153
transform 1 0 6864 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6908
timestamp 1018054153
transform 1 0 6880 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6910
timestamp 1018054153
transform 1 0 6896 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6912
timestamp 1018054153
transform 1 0 6912 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6914
timestamp 1018054153
transform 1 0 6928 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6916
timestamp 1018054153
transform 1 0 6944 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6918
timestamp 1018054153
transform 1 0 6960 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6920
timestamp 1018054153
transform 1 0 6976 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6922
timestamp 1018054153
transform 1 0 6992 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6924
timestamp 1018054153
transform 1 0 7008 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6926
timestamp 1018054153
transform 1 0 7024 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6928
timestamp 1018054153
transform 1 0 7040 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6930
timestamp 1018054153
transform 1 0 7056 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6932
timestamp 1018054153
transform 1 0 7072 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6934
timestamp 1018054153
transform 1 0 7088 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6936
timestamp 1018054153
transform 1 0 7104 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6938
timestamp 1018054153
transform 1 0 7120 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6940
timestamp 1018054153
transform 1 0 7136 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6942
timestamp 1018054153
transform 1 0 7152 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6944
timestamp 1018054153
transform 1 0 7168 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6946
timestamp 1018054153
transform 1 0 7184 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6948
timestamp 1018054153
transform 1 0 7200 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6950
timestamp 1018054153
transform 1 0 7216 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6952
timestamp 1018054153
transform 1 0 7232 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6954
timestamp 1018054153
transform 1 0 7248 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6956
timestamp 1018054153
transform 1 0 7264 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6958
timestamp 1018054153
transform 1 0 7280 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6960
timestamp 1018054153
transform 1 0 7296 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6962
timestamp 1018054153
transform 1 0 7312 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6964
timestamp 1018054153
transform 1 0 7328 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6966
timestamp 1018054153
transform 1 0 7344 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6968
timestamp 1018054153
transform 1 0 7360 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6970
timestamp 1018054153
transform 1 0 7376 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6972
timestamp 1018054153
transform 1 0 7392 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6974
timestamp 1018054153
transform 1 0 7408 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6976
timestamp 1018054153
transform 1 0 7424 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6978
timestamp 1018054153
transform 1 0 7440 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6980
timestamp 1018054153
transform 1 0 7456 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6982
timestamp 1018054153
transform 1 0 7472 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6984
timestamp 1018054153
transform 1 0 7488 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6986
timestamp 1018054153
transform 1 0 7504 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6988
timestamp 1018054153
transform 1 0 7520 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6990
timestamp 1018054153
transform 1 0 7536 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6992
timestamp 1018054153
transform 1 0 7552 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6994
timestamp 1018054153
transform 1 0 7568 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6996
timestamp 1018054153
transform 1 0 7584 0 -1 3280
box -16 -6 32 210
use FILL  FILL_6998
timestamp 1018054153
transform 1 0 7600 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7000
timestamp 1018054153
transform 1 0 7616 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7002
timestamp 1018054153
transform 1 0 7632 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7004
timestamp 1018054153
transform 1 0 7648 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7006
timestamp 1018054153
transform 1 0 7664 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7008
timestamp 1018054153
transform 1 0 7680 0 -1 3280
box -16 -6 32 210
use FILL  FILL_7010
timestamp 1018054153
transform 1 0 7696 0 -1 3280
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_43
timestamp 1542725905
transform 1 0 7788 0 1 3080
box -48 -6 48 6
use FILL  FILL_7012
timestamp 1018054153
transform 1 0 7712 0 -1 3280
box -16 -6 32 210
use M2_M1  M2_M1_288
timestamp 1542725905
transform 1 0 6600 0 1 2930
box -4 -4 4 4
use M2_M1  M2_M1_289
timestamp 1542725905
transform 1 0 7304 0 1 2930
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_44
timestamp 1542725905
transform 1 0 2092 0 1 2880
box -48 -6 48 6
use FILL  FILL_7013
timestamp 1018054153
transform 1 0 2272 0 1 2880
box -16 -6 32 210
use FILL  FILL_7015
timestamp 1018054153
transform 1 0 2288 0 1 2880
box -16 -6 32 210
use FILL  FILL_7017
timestamp 1018054153
transform 1 0 2304 0 1 2880
box -16 -6 32 210
use FILL  FILL_7019
timestamp 1018054153
transform 1 0 2320 0 1 2880
box -16 -6 32 210
use FILL  FILL_7021
timestamp 1018054153
transform 1 0 2336 0 1 2880
box -16 -6 32 210
use FILL  FILL_7023
timestamp 1018054153
transform 1 0 2352 0 1 2880
box -16 -6 32 210
use FILL  FILL_7025
timestamp 1018054153
transform 1 0 2368 0 1 2880
box -16 -6 32 210
use FILL  FILL_7027
timestamp 1018054153
transform 1 0 2384 0 1 2880
box -16 -6 32 210
use FILL  FILL_7029
timestamp 1018054153
transform 1 0 2400 0 1 2880
box -16 -6 32 210
use FILL  FILL_7031
timestamp 1018054153
transform 1 0 2416 0 1 2880
box -16 -6 32 210
use FILL  FILL_7033
timestamp 1018054153
transform 1 0 2432 0 1 2880
box -16 -6 32 210
use FILL  FILL_7035
timestamp 1018054153
transform 1 0 2448 0 1 2880
box -16 -6 32 210
use FILL  FILL_7037
timestamp 1018054153
transform 1 0 2464 0 1 2880
box -16 -6 32 210
use FILL  FILL_7039
timestamp 1018054153
transform 1 0 2480 0 1 2880
box -16 -6 32 210
use FILL  FILL_7041
timestamp 1018054153
transform 1 0 2496 0 1 2880
box -16 -6 32 210
use FILL  FILL_7043
timestamp 1018054153
transform 1 0 2512 0 1 2880
box -16 -6 32 210
use FILL  FILL_7045
timestamp 1018054153
transform 1 0 2528 0 1 2880
box -16 -6 32 210
use FILL  FILL_7047
timestamp 1018054153
transform 1 0 2544 0 1 2880
box -16 -6 32 210
use FILL  FILL_7049
timestamp 1018054153
transform 1 0 2560 0 1 2880
box -16 -6 32 210
use FILL  FILL_7051
timestamp 1018054153
transform 1 0 2576 0 1 2880
box -16 -6 32 210
use FILL  FILL_7053
timestamp 1018054153
transform 1 0 2592 0 1 2880
box -16 -6 32 210
use FILL  FILL_7055
timestamp 1018054153
transform 1 0 2608 0 1 2880
box -16 -6 32 210
use FILL  FILL_7057
timestamp 1018054153
transform 1 0 2624 0 1 2880
box -16 -6 32 210
use FILL  FILL_7059
timestamp 1018054153
transform 1 0 2640 0 1 2880
box -16 -6 32 210
use FILL  FILL_7061
timestamp 1018054153
transform 1 0 2656 0 1 2880
box -16 -6 32 210
use FILL  FILL_7063
timestamp 1018054153
transform 1 0 2672 0 1 2880
box -16 -6 32 210
use FILL  FILL_7065
timestamp 1018054153
transform 1 0 2688 0 1 2880
box -16 -6 32 210
use FILL  FILL_7067
timestamp 1018054153
transform 1 0 2704 0 1 2880
box -16 -6 32 210
use FILL  FILL_7069
timestamp 1018054153
transform 1 0 2720 0 1 2880
box -16 -6 32 210
use FILL  FILL_7071
timestamp 1018054153
transform 1 0 2736 0 1 2880
box -16 -6 32 210
use FILL  FILL_7073
timestamp 1018054153
transform 1 0 2752 0 1 2880
box -16 -6 32 210
use FILL  FILL_7075
timestamp 1018054153
transform 1 0 2768 0 1 2880
box -16 -6 32 210
use FILL  FILL_7077
timestamp 1018054153
transform 1 0 2784 0 1 2880
box -16 -6 32 210
use FILL  FILL_7079
timestamp 1018054153
transform 1 0 2800 0 1 2880
box -16 -6 32 210
use FILL  FILL_7081
timestamp 1018054153
transform 1 0 2816 0 1 2880
box -16 -6 32 210
use FILL  FILL_7083
timestamp 1018054153
transform 1 0 2832 0 1 2880
box -16 -6 32 210
use FILL  FILL_7085
timestamp 1018054153
transform 1 0 2848 0 1 2880
box -16 -6 32 210
use FILL  FILL_7087
timestamp 1018054153
transform 1 0 2864 0 1 2880
box -16 -6 32 210
use FILL  FILL_7089
timestamp 1018054153
transform 1 0 2880 0 1 2880
box -16 -6 32 210
use FILL  FILL_7091
timestamp 1018054153
transform 1 0 2896 0 1 2880
box -16 -6 32 210
use FILL  FILL_7093
timestamp 1018054153
transform 1 0 2912 0 1 2880
box -16 -6 32 210
use FILL  FILL_7095
timestamp 1018054153
transform 1 0 2928 0 1 2880
box -16 -6 32 210
use FILL  FILL_7097
timestamp 1018054153
transform 1 0 2944 0 1 2880
box -16 -6 32 210
use FILL  FILL_7099
timestamp 1018054153
transform 1 0 2960 0 1 2880
box -16 -6 32 210
use FILL  FILL_7101
timestamp 1018054153
transform 1 0 2976 0 1 2880
box -16 -6 32 210
use FILL  FILL_7103
timestamp 1018054153
transform 1 0 2992 0 1 2880
box -16 -6 32 210
use FILL  FILL_7105
timestamp 1018054153
transform 1 0 3008 0 1 2880
box -16 -6 32 210
use FILL  FILL_7107
timestamp 1018054153
transform 1 0 3024 0 1 2880
box -16 -6 32 210
use FILL  FILL_7109
timestamp 1018054153
transform 1 0 3040 0 1 2880
box -16 -6 32 210
use FILL  FILL_7111
timestamp 1018054153
transform 1 0 3056 0 1 2880
box -16 -6 32 210
use FILL  FILL_7113
timestamp 1018054153
transform 1 0 3072 0 1 2880
box -16 -6 32 210
use FILL  FILL_7115
timestamp 1018054153
transform 1 0 3088 0 1 2880
box -16 -6 32 210
use FILL  FILL_7117
timestamp 1018054153
transform 1 0 3104 0 1 2880
box -16 -6 32 210
use FILL  FILL_7119
timestamp 1018054153
transform 1 0 3120 0 1 2880
box -16 -6 32 210
use FILL  FILL_7121
timestamp 1018054153
transform 1 0 3136 0 1 2880
box -16 -6 32 210
use FILL  FILL_7123
timestamp 1018054153
transform 1 0 3152 0 1 2880
box -16 -6 32 210
use FILL  FILL_7125
timestamp 1018054153
transform 1 0 3168 0 1 2880
box -16 -6 32 210
use FILL  FILL_7127
timestamp 1018054153
transform 1 0 3184 0 1 2880
box -16 -6 32 210
use FILL  FILL_7129
timestamp 1018054153
transform 1 0 3200 0 1 2880
box -16 -6 32 210
use FILL  FILL_7131
timestamp 1018054153
transform 1 0 3216 0 1 2880
box -16 -6 32 210
use FILL  FILL_7133
timestamp 1018054153
transform 1 0 3232 0 1 2880
box -16 -6 32 210
use FILL  FILL_7135
timestamp 1018054153
transform 1 0 3248 0 1 2880
box -16 -6 32 210
use FILL  FILL_7137
timestamp 1018054153
transform 1 0 3264 0 1 2880
box -16 -6 32 210
use FILL  FILL_7139
timestamp 1018054153
transform 1 0 3280 0 1 2880
box -16 -6 32 210
use FILL  FILL_7141
timestamp 1018054153
transform 1 0 3296 0 1 2880
box -16 -6 32 210
use FILL  FILL_7143
timestamp 1018054153
transform 1 0 3312 0 1 2880
box -16 -6 32 210
use FILL  FILL_7145
timestamp 1018054153
transform 1 0 3328 0 1 2880
box -16 -6 32 210
use FILL  FILL_7147
timestamp 1018054153
transform 1 0 3344 0 1 2880
box -16 -6 32 210
use FILL  FILL_7149
timestamp 1018054153
transform 1 0 3360 0 1 2880
box -16 -6 32 210
use FILL  FILL_7151
timestamp 1018054153
transform 1 0 3376 0 1 2880
box -16 -6 32 210
use FILL  FILL_7153
timestamp 1018054153
transform 1 0 3392 0 1 2880
box -16 -6 32 210
use FILL  FILL_7155
timestamp 1018054153
transform 1 0 3408 0 1 2880
box -16 -6 32 210
use FILL  FILL_7157
timestamp 1018054153
transform 1 0 3424 0 1 2880
box -16 -6 32 210
use FILL  FILL_7159
timestamp 1018054153
transform 1 0 3440 0 1 2880
box -16 -6 32 210
use FILL  FILL_7161
timestamp 1018054153
transform 1 0 3456 0 1 2880
box -16 -6 32 210
use FILL  FILL_7163
timestamp 1018054153
transform 1 0 3472 0 1 2880
box -16 -6 32 210
use FILL  FILL_7165
timestamp 1018054153
transform 1 0 3488 0 1 2880
box -16 -6 32 210
use FILL  FILL_7167
timestamp 1018054153
transform 1 0 3504 0 1 2880
box -16 -6 32 210
use FILL  FILL_7169
timestamp 1018054153
transform 1 0 3520 0 1 2880
box -16 -6 32 210
use FILL  FILL_7171
timestamp 1018054153
transform 1 0 3536 0 1 2880
box -16 -6 32 210
use FILL  FILL_7173
timestamp 1018054153
transform 1 0 3552 0 1 2880
box -16 -6 32 210
use FILL  FILL_7175
timestamp 1018054153
transform 1 0 3568 0 1 2880
box -16 -6 32 210
use FILL  FILL_7177
timestamp 1018054153
transform 1 0 3584 0 1 2880
box -16 -6 32 210
use FILL  FILL_7179
timestamp 1018054153
transform 1 0 3600 0 1 2880
box -16 -6 32 210
use FILL  FILL_7181
timestamp 1018054153
transform 1 0 3616 0 1 2880
box -16 -6 32 210
use FILL  FILL_7183
timestamp 1018054153
transform 1 0 3632 0 1 2880
box -16 -6 32 210
use FILL  FILL_7185
timestamp 1018054153
transform 1 0 3648 0 1 2880
box -16 -6 32 210
use FILL  FILL_7187
timestamp 1018054153
transform 1 0 3664 0 1 2880
box -16 -6 32 210
use FILL  FILL_7189
timestamp 1018054153
transform 1 0 3680 0 1 2880
box -16 -6 32 210
use FILL  FILL_7191
timestamp 1018054153
transform 1 0 3696 0 1 2880
box -16 -6 32 210
use FILL  FILL_7193
timestamp 1018054153
transform 1 0 3712 0 1 2880
box -16 -6 32 210
use FILL  FILL_7195
timestamp 1018054153
transform 1 0 3728 0 1 2880
box -16 -6 32 210
use FILL  FILL_7197
timestamp 1018054153
transform 1 0 3744 0 1 2880
box -16 -6 32 210
use FILL  FILL_7199
timestamp 1018054153
transform 1 0 3760 0 1 2880
box -16 -6 32 210
use FILL  FILL_7201
timestamp 1018054153
transform 1 0 3776 0 1 2880
box -16 -6 32 210
use FILL  FILL_7203
timestamp 1018054153
transform 1 0 3792 0 1 2880
box -16 -6 32 210
use FILL  FILL_7205
timestamp 1018054153
transform 1 0 3808 0 1 2880
box -16 -6 32 210
use FILL  FILL_7207
timestamp 1018054153
transform 1 0 3824 0 1 2880
box -16 -6 32 210
use FILL  FILL_7209
timestamp 1018054153
transform 1 0 3840 0 1 2880
box -16 -6 32 210
use FILL  FILL_7211
timestamp 1018054153
transform 1 0 3856 0 1 2880
box -16 -6 32 210
use FILL  FILL_7213
timestamp 1018054153
transform 1 0 3872 0 1 2880
box -16 -6 32 210
use FILL  FILL_7215
timestamp 1018054153
transform 1 0 3888 0 1 2880
box -16 -6 32 210
use FILL  FILL_7217
timestamp 1018054153
transform 1 0 3904 0 1 2880
box -16 -6 32 210
use FILL  FILL_7219
timestamp 1018054153
transform 1 0 3920 0 1 2880
box -16 -6 32 210
use FILL  FILL_7221
timestamp 1018054153
transform 1 0 3936 0 1 2880
box -16 -6 32 210
use FILL  FILL_7223
timestamp 1018054153
transform 1 0 3952 0 1 2880
box -16 -6 32 210
use FILL  FILL_7225
timestamp 1018054153
transform 1 0 3968 0 1 2880
box -16 -6 32 210
use FILL  FILL_7227
timestamp 1018054153
transform 1 0 3984 0 1 2880
box -16 -6 32 210
use FILL  FILL_7229
timestamp 1018054153
transform 1 0 4000 0 1 2880
box -16 -6 32 210
use FILL  FILL_7231
timestamp 1018054153
transform 1 0 4016 0 1 2880
box -16 -6 32 210
use FILL  FILL_7233
timestamp 1018054153
transform 1 0 4032 0 1 2880
box -16 -6 32 210
use FILL  FILL_7235
timestamp 1018054153
transform 1 0 4048 0 1 2880
box -16 -6 32 210
use FILL  FILL_7237
timestamp 1018054153
transform 1 0 4064 0 1 2880
box -16 -6 32 210
use FILL  FILL_7239
timestamp 1018054153
transform 1 0 4080 0 1 2880
box -16 -6 32 210
use FILL  FILL_7241
timestamp 1018054153
transform 1 0 4096 0 1 2880
box -16 -6 32 210
use FILL  FILL_7243
timestamp 1018054153
transform 1 0 4112 0 1 2880
box -16 -6 32 210
use FILL  FILL_7245
timestamp 1018054153
transform 1 0 4128 0 1 2880
box -16 -6 32 210
use FILL  FILL_7247
timestamp 1018054153
transform 1 0 4144 0 1 2880
box -16 -6 32 210
use FILL  FILL_7249
timestamp 1018054153
transform 1 0 4160 0 1 2880
box -16 -6 32 210
use FILL  FILL_7251
timestamp 1018054153
transform 1 0 4176 0 1 2880
box -16 -6 32 210
use FILL  FILL_7253
timestamp 1018054153
transform 1 0 4192 0 1 2880
box -16 -6 32 210
use FILL  FILL_7255
timestamp 1018054153
transform 1 0 4208 0 1 2880
box -16 -6 32 210
use FILL  FILL_7257
timestamp 1018054153
transform 1 0 4224 0 1 2880
box -16 -6 32 210
use FILL  FILL_7259
timestamp 1018054153
transform 1 0 4240 0 1 2880
box -16 -6 32 210
use FILL  FILL_7261
timestamp 1018054153
transform 1 0 4256 0 1 2880
box -16 -6 32 210
use FILL  FILL_7263
timestamp 1018054153
transform 1 0 4272 0 1 2880
box -16 -6 32 210
use FILL  FILL_7265
timestamp 1018054153
transform 1 0 4288 0 1 2880
box -16 -6 32 210
use FILL  FILL_7267
timestamp 1018054153
transform 1 0 4304 0 1 2880
box -16 -6 32 210
use FILL  FILL_7269
timestamp 1018054153
transform 1 0 4320 0 1 2880
box -16 -6 32 210
use FILL  FILL_7271
timestamp 1018054153
transform 1 0 4336 0 1 2880
box -16 -6 32 210
use FILL  FILL_7273
timestamp 1018054153
transform 1 0 4352 0 1 2880
box -16 -6 32 210
use FILL  FILL_7275
timestamp 1018054153
transform 1 0 4368 0 1 2880
box -16 -6 32 210
use FILL  FILL_7277
timestamp 1018054153
transform 1 0 4384 0 1 2880
box -16 -6 32 210
use FILL  FILL_7279
timestamp 1018054153
transform 1 0 4400 0 1 2880
box -16 -6 32 210
use FILL  FILL_7281
timestamp 1018054153
transform 1 0 4416 0 1 2880
box -16 -6 32 210
use FILL  FILL_7283
timestamp 1018054153
transform 1 0 4432 0 1 2880
box -16 -6 32 210
use FILL  FILL_7285
timestamp 1018054153
transform 1 0 4448 0 1 2880
box -16 -6 32 210
use FILL  FILL_7287
timestamp 1018054153
transform 1 0 4464 0 1 2880
box -16 -6 32 210
use FILL  FILL_7289
timestamp 1018054153
transform 1 0 4480 0 1 2880
box -16 -6 32 210
use FILL  FILL_7291
timestamp 1018054153
transform 1 0 4496 0 1 2880
box -16 -6 32 210
use FILL  FILL_7293
timestamp 1018054153
transform 1 0 4512 0 1 2880
box -16 -6 32 210
use FILL  FILL_7295
timestamp 1018054153
transform 1 0 4528 0 1 2880
box -16 -6 32 210
use FILL  FILL_7297
timestamp 1018054153
transform 1 0 4544 0 1 2880
box -16 -6 32 210
use FILL  FILL_7299
timestamp 1018054153
transform 1 0 4560 0 1 2880
box -16 -6 32 210
use FILL  FILL_7301
timestamp 1018054153
transform 1 0 4576 0 1 2880
box -16 -6 32 210
use FILL  FILL_7303
timestamp 1018054153
transform 1 0 4592 0 1 2880
box -16 -6 32 210
use FILL  FILL_7305
timestamp 1018054153
transform 1 0 4608 0 1 2880
box -16 -6 32 210
use FILL  FILL_7307
timestamp 1018054153
transform 1 0 4624 0 1 2880
box -16 -6 32 210
use FILL  FILL_7309
timestamp 1018054153
transform 1 0 4640 0 1 2880
box -16 -6 32 210
use FILL  FILL_7311
timestamp 1018054153
transform 1 0 4656 0 1 2880
box -16 -6 32 210
use FILL  FILL_7313
timestamp 1018054153
transform 1 0 4672 0 1 2880
box -16 -6 32 210
use FILL  FILL_7315
timestamp 1018054153
transform 1 0 4688 0 1 2880
box -16 -6 32 210
use FILL  FILL_7317
timestamp 1018054153
transform 1 0 4704 0 1 2880
box -16 -6 32 210
use FILL  FILL_7319
timestamp 1018054153
transform 1 0 4720 0 1 2880
box -16 -6 32 210
use FILL  FILL_7321
timestamp 1018054153
transform 1 0 4736 0 1 2880
box -16 -6 32 210
use FILL  FILL_7323
timestamp 1018054153
transform 1 0 4752 0 1 2880
box -16 -6 32 210
use FILL  FILL_7325
timestamp 1018054153
transform 1 0 4768 0 1 2880
box -16 -6 32 210
use FILL  FILL_7327
timestamp 1018054153
transform 1 0 4784 0 1 2880
box -16 -6 32 210
use FILL  FILL_7329
timestamp 1018054153
transform 1 0 4800 0 1 2880
box -16 -6 32 210
use FILL  FILL_7331
timestamp 1018054153
transform 1 0 4816 0 1 2880
box -16 -6 32 210
use FILL  FILL_7333
timestamp 1018054153
transform 1 0 4832 0 1 2880
box -16 -6 32 210
use FILL  FILL_7335
timestamp 1018054153
transform 1 0 4848 0 1 2880
box -16 -6 32 210
use FILL  FILL_7337
timestamp 1018054153
transform 1 0 4864 0 1 2880
box -16 -6 32 210
use FILL  FILL_7339
timestamp 1018054153
transform 1 0 4880 0 1 2880
box -16 -6 32 210
use FILL  FILL_7341
timestamp 1018054153
transform 1 0 4896 0 1 2880
box -16 -6 32 210
use FILL  FILL_7343
timestamp 1018054153
transform 1 0 4912 0 1 2880
box -16 -6 32 210
use FILL  FILL_7345
timestamp 1018054153
transform 1 0 4928 0 1 2880
box -16 -6 32 210
use FILL  FILL_7347
timestamp 1018054153
transform 1 0 4944 0 1 2880
box -16 -6 32 210
use FILL  FILL_7349
timestamp 1018054153
transform 1 0 4960 0 1 2880
box -16 -6 32 210
use FILL  FILL_7351
timestamp 1018054153
transform 1 0 4976 0 1 2880
box -16 -6 32 210
use FILL  FILL_7353
timestamp 1018054153
transform 1 0 4992 0 1 2880
box -16 -6 32 210
use FILL  FILL_7355
timestamp 1018054153
transform 1 0 5008 0 1 2880
box -16 -6 32 210
use FILL  FILL_7357
timestamp 1018054153
transform 1 0 5024 0 1 2880
box -16 -6 32 210
use FILL  FILL_7359
timestamp 1018054153
transform 1 0 5040 0 1 2880
box -16 -6 32 210
use FILL  FILL_7361
timestamp 1018054153
transform 1 0 5056 0 1 2880
box -16 -6 32 210
use FILL  FILL_7363
timestamp 1018054153
transform 1 0 5072 0 1 2880
box -16 -6 32 210
use FILL  FILL_7365
timestamp 1018054153
transform 1 0 5088 0 1 2880
box -16 -6 32 210
use FILL  FILL_7367
timestamp 1018054153
transform 1 0 5104 0 1 2880
box -16 -6 32 210
use FILL  FILL_7369
timestamp 1018054153
transform 1 0 5120 0 1 2880
box -16 -6 32 210
use FILL  FILL_7371
timestamp 1018054153
transform 1 0 5136 0 1 2880
box -16 -6 32 210
use FILL  FILL_7373
timestamp 1018054153
transform 1 0 5152 0 1 2880
box -16 -6 32 210
use FILL  FILL_7375
timestamp 1018054153
transform 1 0 5168 0 1 2880
box -16 -6 32 210
use FILL  FILL_7377
timestamp 1018054153
transform 1 0 5184 0 1 2880
box -16 -6 32 210
use FILL  FILL_7379
timestamp 1018054153
transform 1 0 5200 0 1 2880
box -16 -6 32 210
use FILL  FILL_7381
timestamp 1018054153
transform 1 0 5216 0 1 2880
box -16 -6 32 210
use FILL  FILL_7383
timestamp 1018054153
transform 1 0 5232 0 1 2880
box -16 -6 32 210
use FILL  FILL_7385
timestamp 1018054153
transform 1 0 5248 0 1 2880
box -16 -6 32 210
use FILL  FILL_7387
timestamp 1018054153
transform 1 0 5264 0 1 2880
box -16 -6 32 210
use FILL  FILL_7389
timestamp 1018054153
transform 1 0 5280 0 1 2880
box -16 -6 32 210
use FILL  FILL_7391
timestamp 1018054153
transform 1 0 5296 0 1 2880
box -16 -6 32 210
use FILL  FILL_7393
timestamp 1018054153
transform 1 0 5312 0 1 2880
box -16 -6 32 210
use FILL  FILL_7395
timestamp 1018054153
transform 1 0 5328 0 1 2880
box -16 -6 32 210
use FILL  FILL_7397
timestamp 1018054153
transform 1 0 5344 0 1 2880
box -16 -6 32 210
use FILL  FILL_7399
timestamp 1018054153
transform 1 0 5360 0 1 2880
box -16 -6 32 210
use FILL  FILL_7401
timestamp 1018054153
transform 1 0 5376 0 1 2880
box -16 -6 32 210
use FILL  FILL_7403
timestamp 1018054153
transform 1 0 5392 0 1 2880
box -16 -6 32 210
use FILL  FILL_7405
timestamp 1018054153
transform 1 0 5408 0 1 2880
box -16 -6 32 210
use FILL  FILL_7407
timestamp 1018054153
transform 1 0 5424 0 1 2880
box -16 -6 32 210
use FILL  FILL_7409
timestamp 1018054153
transform 1 0 5440 0 1 2880
box -16 -6 32 210
use FILL  FILL_7411
timestamp 1018054153
transform 1 0 5456 0 1 2880
box -16 -6 32 210
use FILL  FILL_7413
timestamp 1018054153
transform 1 0 5472 0 1 2880
box -16 -6 32 210
use FILL  FILL_7415
timestamp 1018054153
transform 1 0 5488 0 1 2880
box -16 -6 32 210
use FILL  FILL_7417
timestamp 1018054153
transform 1 0 5504 0 1 2880
box -16 -6 32 210
use FILL  FILL_7419
timestamp 1018054153
transform 1 0 5520 0 1 2880
box -16 -6 32 210
use FILL  FILL_7421
timestamp 1018054153
transform 1 0 5536 0 1 2880
box -16 -6 32 210
use FILL  FILL_7423
timestamp 1018054153
transform 1 0 5552 0 1 2880
box -16 -6 32 210
use FILL  FILL_7425
timestamp 1018054153
transform 1 0 5568 0 1 2880
box -16 -6 32 210
use FILL  FILL_7427
timestamp 1018054153
transform 1 0 5584 0 1 2880
box -16 -6 32 210
use FILL  FILL_7429
timestamp 1018054153
transform 1 0 5600 0 1 2880
box -16 -6 32 210
use FILL  FILL_7431
timestamp 1018054153
transform 1 0 5616 0 1 2880
box -16 -6 32 210
use FILL  FILL_7433
timestamp 1018054153
transform 1 0 5632 0 1 2880
box -16 -6 32 210
use FILL  FILL_7435
timestamp 1018054153
transform 1 0 5648 0 1 2880
box -16 -6 32 210
use FILL  FILL_7437
timestamp 1018054153
transform 1 0 5664 0 1 2880
box -16 -6 32 210
use FILL  FILL_7439
timestamp 1018054153
transform 1 0 5680 0 1 2880
box -16 -6 32 210
use FILL  FILL_7441
timestamp 1018054153
transform 1 0 5696 0 1 2880
box -16 -6 32 210
use FILL  FILL_7443
timestamp 1018054153
transform 1 0 5712 0 1 2880
box -16 -6 32 210
use FILL  FILL_7445
timestamp 1018054153
transform 1 0 5728 0 1 2880
box -16 -6 32 210
use FILL  FILL_7447
timestamp 1018054153
transform 1 0 5744 0 1 2880
box -16 -6 32 210
use FILL  FILL_7449
timestamp 1018054153
transform 1 0 5760 0 1 2880
box -16 -6 32 210
use FILL  FILL_7451
timestamp 1018054153
transform 1 0 5776 0 1 2880
box -16 -6 32 210
use FILL  FILL_7453
timestamp 1018054153
transform 1 0 5792 0 1 2880
box -16 -6 32 210
use FILL  FILL_7455
timestamp 1018054153
transform 1 0 5808 0 1 2880
box -16 -6 32 210
use FILL  FILL_7457
timestamp 1018054153
transform 1 0 5824 0 1 2880
box -16 -6 32 210
use FILL  FILL_7459
timestamp 1018054153
transform 1 0 5840 0 1 2880
box -16 -6 32 210
use FILL  FILL_7461
timestamp 1018054153
transform 1 0 5856 0 1 2880
box -16 -6 32 210
use FILL  FILL_7463
timestamp 1018054153
transform 1 0 5872 0 1 2880
box -16 -6 32 210
use FILL  FILL_7465
timestamp 1018054153
transform 1 0 5888 0 1 2880
box -16 -6 32 210
use FILL  FILL_7467
timestamp 1018054153
transform 1 0 5904 0 1 2880
box -16 -6 32 210
use FILL  FILL_7469
timestamp 1018054153
transform 1 0 5920 0 1 2880
box -16 -6 32 210
use FILL  FILL_7471
timestamp 1018054153
transform 1 0 5936 0 1 2880
box -16 -6 32 210
use FILL  FILL_7473
timestamp 1018054153
transform 1 0 5952 0 1 2880
box -16 -6 32 210
use FILL  FILL_7475
timestamp 1018054153
transform 1 0 5968 0 1 2880
box -16 -6 32 210
use FILL  FILL_7477
timestamp 1018054153
transform 1 0 5984 0 1 2880
box -16 -6 32 210
use FILL  FILL_7479
timestamp 1018054153
transform 1 0 6000 0 1 2880
box -16 -6 32 210
use FILL  FILL_7481
timestamp 1018054153
transform 1 0 6016 0 1 2880
box -16 -6 32 210
use FILL  FILL_7483
timestamp 1018054153
transform 1 0 6032 0 1 2880
box -16 -6 32 210
use FILL  FILL_7485
timestamp 1018054153
transform 1 0 6048 0 1 2880
box -16 -6 32 210
use FILL  FILL_7487
timestamp 1018054153
transform 1 0 6064 0 1 2880
box -16 -6 32 210
use FILL  FILL_7489
timestamp 1018054153
transform 1 0 6080 0 1 2880
box -16 -6 32 210
use FILL  FILL_7491
timestamp 1018054153
transform 1 0 6096 0 1 2880
box -16 -6 32 210
use FILL  FILL_7493
timestamp 1018054153
transform 1 0 6112 0 1 2880
box -16 -6 32 210
use FILL  FILL_7495
timestamp 1018054153
transform 1 0 6128 0 1 2880
box -16 -6 32 210
use FILL  FILL_7497
timestamp 1018054153
transform 1 0 6144 0 1 2880
box -16 -6 32 210
use FILL  FILL_7499
timestamp 1018054153
transform 1 0 6160 0 1 2880
box -16 -6 32 210
use FILL  FILL_7501
timestamp 1018054153
transform 1 0 6176 0 1 2880
box -16 -6 32 210
use FILL  FILL_7503
timestamp 1018054153
transform 1 0 6192 0 1 2880
box -16 -6 32 210
use FILL  FILL_7505
timestamp 1018054153
transform 1 0 6208 0 1 2880
box -16 -6 32 210
use FILL  FILL_7507
timestamp 1018054153
transform 1 0 6224 0 1 2880
box -16 -6 32 210
use FILL  FILL_7509
timestamp 1018054153
transform 1 0 6240 0 1 2880
box -16 -6 32 210
use FILL  FILL_7511
timestamp 1018054153
transform 1 0 6256 0 1 2880
box -16 -6 32 210
use FILL  FILL_7513
timestamp 1018054153
transform 1 0 6272 0 1 2880
box -16 -6 32 210
use FILL  FILL_7515
timestamp 1018054153
transform 1 0 6288 0 1 2880
box -16 -6 32 210
use FILL  FILL_7517
timestamp 1018054153
transform 1 0 6304 0 1 2880
box -16 -6 32 210
use FILL  FILL_7519
timestamp 1018054153
transform 1 0 6320 0 1 2880
box -16 -6 32 210
use FILL  FILL_7521
timestamp 1018054153
transform 1 0 6336 0 1 2880
box -16 -6 32 210
use FILL  FILL_7523
timestamp 1018054153
transform 1 0 6352 0 1 2880
box -16 -6 32 210
use FILL  FILL_7525
timestamp 1018054153
transform 1 0 6368 0 1 2880
box -16 -6 32 210
use FILL  FILL_7527
timestamp 1018054153
transform 1 0 6384 0 1 2880
box -16 -6 32 210
use FILL  FILL_7529
timestamp 1018054153
transform 1 0 6400 0 1 2880
box -16 -6 32 210
use FILL  FILL_7531
timestamp 1018054153
transform 1 0 6416 0 1 2880
box -16 -6 32 210
use FILL  FILL_7533
timestamp 1018054153
transform 1 0 6432 0 1 2880
box -16 -6 32 210
use FILL  FILL_7535
timestamp 1018054153
transform 1 0 6448 0 1 2880
box -16 -6 32 210
use FILL  FILL_7537
timestamp 1018054153
transform 1 0 6464 0 1 2880
box -16 -6 32 210
use FILL  FILL_7539
timestamp 1018054153
transform 1 0 6480 0 1 2880
box -16 -6 32 210
use FILL  FILL_7541
timestamp 1018054153
transform 1 0 6496 0 1 2880
box -16 -6 32 210
use FILL  FILL_7543
timestamp 1018054153
transform 1 0 6512 0 1 2880
box -16 -6 32 210
use FILL  FILL_7545
timestamp 1018054153
transform 1 0 6528 0 1 2880
box -16 -6 32 210
use FILL  FILL_7547
timestamp 1018054153
transform 1 0 6544 0 1 2880
box -16 -6 32 210
use FILL  FILL_7549
timestamp 1018054153
transform 1 0 6560 0 1 2880
box -16 -6 32 210
use FILL  FILL_7551
timestamp 1018054153
transform 1 0 6576 0 1 2880
box -16 -6 32 210
use FILL  FILL_7553
timestamp 1018054153
transform 1 0 6592 0 1 2880
box -16 -6 32 210
use FILL  FILL_7555
timestamp 1018054153
transform 1 0 6608 0 1 2880
box -16 -6 32 210
use FILL  FILL_7557
timestamp 1018054153
transform 1 0 6624 0 1 2880
box -16 -6 32 210
use FILL  FILL_7559
timestamp 1018054153
transform 1 0 6640 0 1 2880
box -16 -6 32 210
use FILL  FILL_7561
timestamp 1018054153
transform 1 0 6656 0 1 2880
box -16 -6 32 210
use FILL  FILL_7563
timestamp 1018054153
transform 1 0 6672 0 1 2880
box -16 -6 32 210
use FILL  FILL_7565
timestamp 1018054153
transform 1 0 6688 0 1 2880
box -16 -6 32 210
use FILL  FILL_7567
timestamp 1018054153
transform 1 0 6704 0 1 2880
box -16 -6 32 210
use FILL  FILL_7569
timestamp 1018054153
transform 1 0 6720 0 1 2880
box -16 -6 32 210
use FILL  FILL_7571
timestamp 1018054153
transform 1 0 6736 0 1 2880
box -16 -6 32 210
use FILL  FILL_7573
timestamp 1018054153
transform 1 0 6752 0 1 2880
box -16 -6 32 210
use FILL  FILL_7575
timestamp 1018054153
transform 1 0 6768 0 1 2880
box -16 -6 32 210
use FILL  FILL_7577
timestamp 1018054153
transform 1 0 6784 0 1 2880
box -16 -6 32 210
use FILL  FILL_7579
timestamp 1018054153
transform 1 0 6800 0 1 2880
box -16 -6 32 210
use FILL  FILL_7581
timestamp 1018054153
transform 1 0 6816 0 1 2880
box -16 -6 32 210
use FILL  FILL_7583
timestamp 1018054153
transform 1 0 6832 0 1 2880
box -16 -6 32 210
use FILL  FILL_7585
timestamp 1018054153
transform 1 0 6848 0 1 2880
box -16 -6 32 210
use FILL  FILL_7587
timestamp 1018054153
transform 1 0 6864 0 1 2880
box -16 -6 32 210
use FILL  FILL_7589
timestamp 1018054153
transform 1 0 6880 0 1 2880
box -16 -6 32 210
use FILL  FILL_7591
timestamp 1018054153
transform 1 0 6896 0 1 2880
box -16 -6 32 210
use FILL  FILL_7593
timestamp 1018054153
transform 1 0 6912 0 1 2880
box -16 -6 32 210
use FILL  FILL_7595
timestamp 1018054153
transform 1 0 6928 0 1 2880
box -16 -6 32 210
use FILL  FILL_7597
timestamp 1018054153
transform 1 0 6944 0 1 2880
box -16 -6 32 210
use FILL  FILL_7599
timestamp 1018054153
transform 1 0 6960 0 1 2880
box -16 -6 32 210
use FILL  FILL_7601
timestamp 1018054153
transform 1 0 6976 0 1 2880
box -16 -6 32 210
use FILL  FILL_7603
timestamp 1018054153
transform 1 0 6992 0 1 2880
box -16 -6 32 210
use FILL  FILL_7605
timestamp 1018054153
transform 1 0 7008 0 1 2880
box -16 -6 32 210
use FILL  FILL_7607
timestamp 1018054153
transform 1 0 7024 0 1 2880
box -16 -6 32 210
use FILL  FILL_7609
timestamp 1018054153
transform 1 0 7040 0 1 2880
box -16 -6 32 210
use FILL  FILL_7611
timestamp 1018054153
transform 1 0 7056 0 1 2880
box -16 -6 32 210
use FILL  FILL_7613
timestamp 1018054153
transform 1 0 7072 0 1 2880
box -16 -6 32 210
use FILL  FILL_7615
timestamp 1018054153
transform 1 0 7088 0 1 2880
box -16 -6 32 210
use FILL  FILL_7617
timestamp 1018054153
transform 1 0 7104 0 1 2880
box -16 -6 32 210
use FILL  FILL_7619
timestamp 1018054153
transform 1 0 7120 0 1 2880
box -16 -6 32 210
use FILL  FILL_7621
timestamp 1018054153
transform 1 0 7136 0 1 2880
box -16 -6 32 210
use FILL  FILL_7623
timestamp 1018054153
transform 1 0 7152 0 1 2880
box -16 -6 32 210
use FILL  FILL_7625
timestamp 1018054153
transform 1 0 7168 0 1 2880
box -16 -6 32 210
use FILL  FILL_7627
timestamp 1018054153
transform 1 0 7184 0 1 2880
box -16 -6 32 210
use FILL  FILL_7629
timestamp 1018054153
transform 1 0 7200 0 1 2880
box -16 -6 32 210
use FILL  FILL_7631
timestamp 1018054153
transform 1 0 7216 0 1 2880
box -16 -6 32 210
use FILL  FILL_7633
timestamp 1018054153
transform 1 0 7232 0 1 2880
box -16 -6 32 210
use FILL  FILL_7635
timestamp 1018054153
transform 1 0 7248 0 1 2880
box -16 -6 32 210
use FILL  FILL_7637
timestamp 1018054153
transform 1 0 7264 0 1 2880
box -16 -6 32 210
use FILL  FILL_7639
timestamp 1018054153
transform 1 0 7280 0 1 2880
box -16 -6 32 210
use FILL  FILL_7641
timestamp 1018054153
transform 1 0 7296 0 1 2880
box -16 -6 32 210
use FILL  FILL_7643
timestamp 1018054153
transform 1 0 7312 0 1 2880
box -16 -6 32 210
use FILL  FILL_7645
timestamp 1018054153
transform 1 0 7328 0 1 2880
box -16 -6 32 210
use FILL  FILL_7647
timestamp 1018054153
transform 1 0 7344 0 1 2880
box -16 -6 32 210
use FILL  FILL_7649
timestamp 1018054153
transform 1 0 7360 0 1 2880
box -16 -6 32 210
use FILL  FILL_7651
timestamp 1018054153
transform 1 0 7376 0 1 2880
box -16 -6 32 210
use FILL  FILL_7653
timestamp 1018054153
transform 1 0 7392 0 1 2880
box -16 -6 32 210
use FILL  FILL_7655
timestamp 1018054153
transform 1 0 7408 0 1 2880
box -16 -6 32 210
use FILL  FILL_7657
timestamp 1018054153
transform 1 0 7424 0 1 2880
box -16 -6 32 210
use FILL  FILL_7659
timestamp 1018054153
transform 1 0 7440 0 1 2880
box -16 -6 32 210
use FILL  FILL_7661
timestamp 1018054153
transform 1 0 7456 0 1 2880
box -16 -6 32 210
use FILL  FILL_7663
timestamp 1018054153
transform 1 0 7472 0 1 2880
box -16 -6 32 210
use FILL  FILL_7665
timestamp 1018054153
transform 1 0 7488 0 1 2880
box -16 -6 32 210
use FILL  FILL_7667
timestamp 1018054153
transform 1 0 7504 0 1 2880
box -16 -6 32 210
use FILL  FILL_7669
timestamp 1018054153
transform 1 0 7520 0 1 2880
box -16 -6 32 210
use FILL  FILL_7671
timestamp 1018054153
transform 1 0 7536 0 1 2880
box -16 -6 32 210
use FILL  FILL_7673
timestamp 1018054153
transform 1 0 7552 0 1 2880
box -16 -6 32 210
use FILL  FILL_7675
timestamp 1018054153
transform 1 0 7568 0 1 2880
box -16 -6 32 210
use FILL  FILL_7677
timestamp 1018054153
transform 1 0 7584 0 1 2880
box -16 -6 32 210
use FILL  FILL_7679
timestamp 1018054153
transform 1 0 7600 0 1 2880
box -16 -6 32 210
use FILL  FILL_7681
timestamp 1018054153
transform 1 0 7616 0 1 2880
box -16 -6 32 210
use FILL  FILL_7683
timestamp 1018054153
transform 1 0 7632 0 1 2880
box -16 -6 32 210
use FILL  FILL_7685
timestamp 1018054153
transform 1 0 7648 0 1 2880
box -16 -6 32 210
use FILL  FILL_7687
timestamp 1018054153
transform 1 0 7664 0 1 2880
box -16 -6 32 210
use FILL  FILL_7689
timestamp 1018054153
transform 1 0 7680 0 1 2880
box -16 -6 32 210
use FILL  FILL_7691
timestamp 1018054153
transform 1 0 7696 0 1 2880
box -16 -6 32 210
use FILL  FILL_7693
timestamp 1018054153
transform 1 0 7712 0 1 2880
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_45
timestamp 1542725905
transform 1 0 7908 0 1 2880
box -48 -6 48 6
use mult_pad_VIA1  mult_pad_VIA1_46
timestamp 1542725905
transform 1 0 2212 0 1 2680
box -48 -6 48 6
use PADNC  PADNC_8
timestamp 1084294400
transform 0 -1 2000 1 0 2600
box -6 -6 606 2000
use FILL  FILL_7014
timestamp 1018054153
transform 1 0 2272 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7016
timestamp 1018054153
transform 1 0 2288 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7018
timestamp 1018054153
transform 1 0 2304 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7020
timestamp 1018054153
transform 1 0 2320 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7022
timestamp 1018054153
transform 1 0 2336 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7024
timestamp 1018054153
transform 1 0 2352 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7026
timestamp 1018054153
transform 1 0 2368 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7028
timestamp 1018054153
transform 1 0 2384 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7030
timestamp 1018054153
transform 1 0 2400 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7032
timestamp 1018054153
transform 1 0 2416 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7034
timestamp 1018054153
transform 1 0 2432 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7036
timestamp 1018054153
transform 1 0 2448 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7038
timestamp 1018054153
transform 1 0 2464 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7040
timestamp 1018054153
transform 1 0 2480 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7042
timestamp 1018054153
transform 1 0 2496 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7044
timestamp 1018054153
transform 1 0 2512 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7046
timestamp 1018054153
transform 1 0 2528 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7048
timestamp 1018054153
transform 1 0 2544 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7050
timestamp 1018054153
transform 1 0 2560 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7052
timestamp 1018054153
transform 1 0 2576 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7054
timestamp 1018054153
transform 1 0 2592 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7056
timestamp 1018054153
transform 1 0 2608 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7058
timestamp 1018054153
transform 1 0 2624 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7060
timestamp 1018054153
transform 1 0 2640 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7062
timestamp 1018054153
transform 1 0 2656 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7064
timestamp 1018054153
transform 1 0 2672 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7066
timestamp 1018054153
transform 1 0 2688 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7068
timestamp 1018054153
transform 1 0 2704 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7070
timestamp 1018054153
transform 1 0 2720 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7072
timestamp 1018054153
transform 1 0 2736 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7074
timestamp 1018054153
transform 1 0 2752 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7076
timestamp 1018054153
transform 1 0 2768 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7078
timestamp 1018054153
transform 1 0 2784 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7080
timestamp 1018054153
transform 1 0 2800 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7082
timestamp 1018054153
transform 1 0 2816 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7084
timestamp 1018054153
transform 1 0 2832 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7086
timestamp 1018054153
transform 1 0 2848 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7088
timestamp 1018054153
transform 1 0 2864 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7090
timestamp 1018054153
transform 1 0 2880 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7092
timestamp 1018054153
transform 1 0 2896 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7094
timestamp 1018054153
transform 1 0 2912 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7096
timestamp 1018054153
transform 1 0 2928 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7098
timestamp 1018054153
transform 1 0 2944 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7100
timestamp 1018054153
transform 1 0 2960 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7102
timestamp 1018054153
transform 1 0 2976 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7104
timestamp 1018054153
transform 1 0 2992 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7106
timestamp 1018054153
transform 1 0 3008 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7108
timestamp 1018054153
transform 1 0 3024 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7110
timestamp 1018054153
transform 1 0 3040 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7112
timestamp 1018054153
transform 1 0 3056 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7114
timestamp 1018054153
transform 1 0 3072 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7116
timestamp 1018054153
transform 1 0 3088 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7118
timestamp 1018054153
transform 1 0 3104 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7120
timestamp 1018054153
transform 1 0 3120 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7122
timestamp 1018054153
transform 1 0 3136 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7124
timestamp 1018054153
transform 1 0 3152 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7126
timestamp 1018054153
transform 1 0 3168 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7128
timestamp 1018054153
transform 1 0 3184 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7130
timestamp 1018054153
transform 1 0 3200 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7132
timestamp 1018054153
transform 1 0 3216 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7134
timestamp 1018054153
transform 1 0 3232 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7136
timestamp 1018054153
transform 1 0 3248 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7138
timestamp 1018054153
transform 1 0 3264 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7140
timestamp 1018054153
transform 1 0 3280 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7142
timestamp 1018054153
transform 1 0 3296 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7144
timestamp 1018054153
transform 1 0 3312 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7146
timestamp 1018054153
transform 1 0 3328 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7148
timestamp 1018054153
transform 1 0 3344 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7150
timestamp 1018054153
transform 1 0 3360 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7152
timestamp 1018054153
transform 1 0 3376 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7154
timestamp 1018054153
transform 1 0 3392 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7156
timestamp 1018054153
transform 1 0 3408 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7158
timestamp 1018054153
transform 1 0 3424 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7160
timestamp 1018054153
transform 1 0 3440 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7162
timestamp 1018054153
transform 1 0 3456 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7164
timestamp 1018054153
transform 1 0 3472 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7166
timestamp 1018054153
transform 1 0 3488 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7168
timestamp 1018054153
transform 1 0 3504 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7170
timestamp 1018054153
transform 1 0 3520 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7172
timestamp 1018054153
transform 1 0 3536 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7174
timestamp 1018054153
transform 1 0 3552 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7176
timestamp 1018054153
transform 1 0 3568 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7178
timestamp 1018054153
transform 1 0 3584 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7180
timestamp 1018054153
transform 1 0 3600 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7182
timestamp 1018054153
transform 1 0 3616 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7184
timestamp 1018054153
transform 1 0 3632 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7186
timestamp 1018054153
transform 1 0 3648 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7188
timestamp 1018054153
transform 1 0 3664 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7190
timestamp 1018054153
transform 1 0 3680 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7192
timestamp 1018054153
transform 1 0 3696 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7194
timestamp 1018054153
transform 1 0 3712 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7196
timestamp 1018054153
transform 1 0 3728 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7198
timestamp 1018054153
transform 1 0 3744 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7200
timestamp 1018054153
transform 1 0 3760 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7202
timestamp 1018054153
transform 1 0 3776 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7204
timestamp 1018054153
transform 1 0 3792 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7206
timestamp 1018054153
transform 1 0 3808 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7208
timestamp 1018054153
transform 1 0 3824 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7210
timestamp 1018054153
transform 1 0 3840 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7212
timestamp 1018054153
transform 1 0 3856 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7214
timestamp 1018054153
transform 1 0 3872 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7216
timestamp 1018054153
transform 1 0 3888 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7218
timestamp 1018054153
transform 1 0 3904 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7220
timestamp 1018054153
transform 1 0 3920 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7222
timestamp 1018054153
transform 1 0 3936 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7224
timestamp 1018054153
transform 1 0 3952 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7226
timestamp 1018054153
transform 1 0 3968 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7228
timestamp 1018054153
transform 1 0 3984 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7230
timestamp 1018054153
transform 1 0 4000 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7232
timestamp 1018054153
transform 1 0 4016 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7234
timestamp 1018054153
transform 1 0 4032 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7236
timestamp 1018054153
transform 1 0 4048 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7238
timestamp 1018054153
transform 1 0 4064 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7240
timestamp 1018054153
transform 1 0 4080 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7242
timestamp 1018054153
transform 1 0 4096 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7244
timestamp 1018054153
transform 1 0 4112 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7246
timestamp 1018054153
transform 1 0 4128 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7248
timestamp 1018054153
transform 1 0 4144 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7250
timestamp 1018054153
transform 1 0 4160 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7252
timestamp 1018054153
transform 1 0 4176 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7254
timestamp 1018054153
transform 1 0 4192 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7256
timestamp 1018054153
transform 1 0 4208 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7258
timestamp 1018054153
transform 1 0 4224 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7260
timestamp 1018054153
transform 1 0 4240 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7262
timestamp 1018054153
transform 1 0 4256 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7264
timestamp 1018054153
transform 1 0 4272 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7266
timestamp 1018054153
transform 1 0 4288 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7268
timestamp 1018054153
transform 1 0 4304 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7270
timestamp 1018054153
transform 1 0 4320 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7272
timestamp 1018054153
transform 1 0 4336 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7274
timestamp 1018054153
transform 1 0 4352 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7276
timestamp 1018054153
transform 1 0 4368 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7278
timestamp 1018054153
transform 1 0 4384 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7280
timestamp 1018054153
transform 1 0 4400 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7282
timestamp 1018054153
transform 1 0 4416 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7284
timestamp 1018054153
transform 1 0 4432 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7286
timestamp 1018054153
transform 1 0 4448 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7288
timestamp 1018054153
transform 1 0 4464 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7290
timestamp 1018054153
transform 1 0 4480 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7292
timestamp 1018054153
transform 1 0 4496 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7294
timestamp 1018054153
transform 1 0 4512 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7296
timestamp 1018054153
transform 1 0 4528 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7298
timestamp 1018054153
transform 1 0 4544 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7300
timestamp 1018054153
transform 1 0 4560 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7302
timestamp 1018054153
transform 1 0 4576 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7304
timestamp 1018054153
transform 1 0 4592 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7306
timestamp 1018054153
transform 1 0 4608 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7308
timestamp 1018054153
transform 1 0 4624 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7310
timestamp 1018054153
transform 1 0 4640 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7312
timestamp 1018054153
transform 1 0 4656 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7314
timestamp 1018054153
transform 1 0 4672 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7316
timestamp 1018054153
transform 1 0 4688 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7318
timestamp 1018054153
transform 1 0 4704 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7320
timestamp 1018054153
transform 1 0 4720 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7322
timestamp 1018054153
transform 1 0 4736 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7324
timestamp 1018054153
transform 1 0 4752 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7326
timestamp 1018054153
transform 1 0 4768 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7328
timestamp 1018054153
transform 1 0 4784 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7330
timestamp 1018054153
transform 1 0 4800 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7332
timestamp 1018054153
transform 1 0 4816 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7334
timestamp 1018054153
transform 1 0 4832 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7336
timestamp 1018054153
transform 1 0 4848 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7338
timestamp 1018054153
transform 1 0 4864 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7340
timestamp 1018054153
transform 1 0 4880 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7342
timestamp 1018054153
transform 1 0 4896 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7344
timestamp 1018054153
transform 1 0 4912 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7346
timestamp 1018054153
transform 1 0 4928 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7348
timestamp 1018054153
transform 1 0 4944 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7350
timestamp 1018054153
transform 1 0 4960 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7352
timestamp 1018054153
transform 1 0 4976 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7354
timestamp 1018054153
transform 1 0 4992 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7356
timestamp 1018054153
transform 1 0 5008 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7358
timestamp 1018054153
transform 1 0 5024 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7360
timestamp 1018054153
transform 1 0 5040 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7362
timestamp 1018054153
transform 1 0 5056 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7364
timestamp 1018054153
transform 1 0 5072 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7366
timestamp 1018054153
transform 1 0 5088 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7368
timestamp 1018054153
transform 1 0 5104 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7370
timestamp 1018054153
transform 1 0 5120 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7372
timestamp 1018054153
transform 1 0 5136 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7374
timestamp 1018054153
transform 1 0 5152 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7376
timestamp 1018054153
transform 1 0 5168 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7378
timestamp 1018054153
transform 1 0 5184 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7380
timestamp 1018054153
transform 1 0 5200 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7382
timestamp 1018054153
transform 1 0 5216 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7384
timestamp 1018054153
transform 1 0 5232 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7386
timestamp 1018054153
transform 1 0 5248 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7388
timestamp 1018054153
transform 1 0 5264 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7390
timestamp 1018054153
transform 1 0 5280 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7392
timestamp 1018054153
transform 1 0 5296 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7394
timestamp 1018054153
transform 1 0 5312 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7396
timestamp 1018054153
transform 1 0 5328 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7398
timestamp 1018054153
transform 1 0 5344 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7400
timestamp 1018054153
transform 1 0 5360 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7402
timestamp 1018054153
transform 1 0 5376 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7404
timestamp 1018054153
transform 1 0 5392 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7406
timestamp 1018054153
transform 1 0 5408 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7408
timestamp 1018054153
transform 1 0 5424 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7410
timestamp 1018054153
transform 1 0 5440 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7412
timestamp 1018054153
transform 1 0 5456 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7414
timestamp 1018054153
transform 1 0 5472 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7416
timestamp 1018054153
transform 1 0 5488 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7418
timestamp 1018054153
transform 1 0 5504 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7420
timestamp 1018054153
transform 1 0 5520 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7422
timestamp 1018054153
transform 1 0 5536 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7424
timestamp 1018054153
transform 1 0 5552 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7426
timestamp 1018054153
transform 1 0 5568 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7428
timestamp 1018054153
transform 1 0 5584 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7430
timestamp 1018054153
transform 1 0 5600 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7432
timestamp 1018054153
transform 1 0 5616 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7434
timestamp 1018054153
transform 1 0 5632 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7436
timestamp 1018054153
transform 1 0 5648 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7438
timestamp 1018054153
transform 1 0 5664 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7440
timestamp 1018054153
transform 1 0 5680 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7442
timestamp 1018054153
transform 1 0 5696 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7444
timestamp 1018054153
transform 1 0 5712 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7446
timestamp 1018054153
transform 1 0 5728 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7448
timestamp 1018054153
transform 1 0 5744 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7450
timestamp 1018054153
transform 1 0 5760 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7452
timestamp 1018054153
transform 1 0 5776 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7454
timestamp 1018054153
transform 1 0 5792 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7456
timestamp 1018054153
transform 1 0 5808 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7458
timestamp 1018054153
transform 1 0 5824 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7460
timestamp 1018054153
transform 1 0 5840 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7462
timestamp 1018054153
transform 1 0 5856 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7464
timestamp 1018054153
transform 1 0 5872 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7466
timestamp 1018054153
transform 1 0 5888 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7468
timestamp 1018054153
transform 1 0 5904 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7470
timestamp 1018054153
transform 1 0 5920 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7472
timestamp 1018054153
transform 1 0 5936 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7474
timestamp 1018054153
transform 1 0 5952 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7476
timestamp 1018054153
transform 1 0 5968 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7478
timestamp 1018054153
transform 1 0 5984 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7480
timestamp 1018054153
transform 1 0 6000 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7482
timestamp 1018054153
transform 1 0 6016 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7484
timestamp 1018054153
transform 1 0 6032 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7486
timestamp 1018054153
transform 1 0 6048 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7488
timestamp 1018054153
transform 1 0 6064 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7490
timestamp 1018054153
transform 1 0 6080 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7492
timestamp 1018054153
transform 1 0 6096 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7494
timestamp 1018054153
transform 1 0 6112 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7496
timestamp 1018054153
transform 1 0 6128 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7498
timestamp 1018054153
transform 1 0 6144 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7500
timestamp 1018054153
transform 1 0 6160 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7502
timestamp 1018054153
transform 1 0 6176 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7504
timestamp 1018054153
transform 1 0 6192 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7506
timestamp 1018054153
transform 1 0 6208 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7508
timestamp 1018054153
transform 1 0 6224 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7510
timestamp 1018054153
transform 1 0 6240 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7512
timestamp 1018054153
transform 1 0 6256 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7514
timestamp 1018054153
transform 1 0 6272 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7516
timestamp 1018054153
transform 1 0 6288 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7518
timestamp 1018054153
transform 1 0 6304 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7520
timestamp 1018054153
transform 1 0 6320 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7522
timestamp 1018054153
transform 1 0 6336 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7524
timestamp 1018054153
transform 1 0 6352 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7526
timestamp 1018054153
transform 1 0 6368 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7528
timestamp 1018054153
transform 1 0 6384 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7530
timestamp 1018054153
transform 1 0 6400 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7532
timestamp 1018054153
transform 1 0 6416 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7534
timestamp 1018054153
transform 1 0 6432 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7536
timestamp 1018054153
transform 1 0 6448 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7538
timestamp 1018054153
transform 1 0 6464 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7540
timestamp 1018054153
transform 1 0 6480 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7542
timestamp 1018054153
transform 1 0 6496 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7544
timestamp 1018054153
transform 1 0 6512 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7546
timestamp 1018054153
transform 1 0 6528 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7548
timestamp 1018054153
transform 1 0 6544 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7550
timestamp 1018054153
transform 1 0 6560 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7552
timestamp 1018054153
transform 1 0 6576 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7554
timestamp 1018054153
transform 1 0 6592 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7556
timestamp 1018054153
transform 1 0 6608 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7558
timestamp 1018054153
transform 1 0 6624 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7560
timestamp 1018054153
transform 1 0 6640 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7562
timestamp 1018054153
transform 1 0 6656 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7564
timestamp 1018054153
transform 1 0 6672 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7566
timestamp 1018054153
transform 1 0 6688 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7568
timestamp 1018054153
transform 1 0 6704 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7570
timestamp 1018054153
transform 1 0 6720 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7572
timestamp 1018054153
transform 1 0 6736 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7574
timestamp 1018054153
transform 1 0 6752 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7576
timestamp 1018054153
transform 1 0 6768 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7578
timestamp 1018054153
transform 1 0 6784 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7580
timestamp 1018054153
transform 1 0 6800 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7582
timestamp 1018054153
transform 1 0 6816 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7584
timestamp 1018054153
transform 1 0 6832 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7586
timestamp 1018054153
transform 1 0 6848 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7588
timestamp 1018054153
transform 1 0 6864 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7590
timestamp 1018054153
transform 1 0 6880 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7592
timestamp 1018054153
transform 1 0 6896 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7594
timestamp 1018054153
transform 1 0 6912 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7596
timestamp 1018054153
transform 1 0 6928 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7598
timestamp 1018054153
transform 1 0 6944 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7600
timestamp 1018054153
transform 1 0 6960 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7602
timestamp 1018054153
transform 1 0 6976 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7604
timestamp 1018054153
transform 1 0 6992 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7606
timestamp 1018054153
transform 1 0 7008 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7608
timestamp 1018054153
transform 1 0 7024 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7610
timestamp 1018054153
transform 1 0 7040 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7612
timestamp 1018054153
transform 1 0 7056 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7614
timestamp 1018054153
transform 1 0 7072 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7616
timestamp 1018054153
transform 1 0 7088 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7618
timestamp 1018054153
transform 1 0 7104 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7620
timestamp 1018054153
transform 1 0 7120 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7622
timestamp 1018054153
transform 1 0 7136 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7624
timestamp 1018054153
transform 1 0 7152 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7626
timestamp 1018054153
transform 1 0 7168 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7628
timestamp 1018054153
transform 1 0 7184 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7630
timestamp 1018054153
transform 1 0 7200 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7632
timestamp 1018054153
transform 1 0 7216 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7634
timestamp 1018054153
transform 1 0 7232 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7636
timestamp 1018054153
transform 1 0 7248 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7638
timestamp 1018054153
transform 1 0 7264 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7640
timestamp 1018054153
transform 1 0 7280 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7642
timestamp 1018054153
transform 1 0 7296 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7644
timestamp 1018054153
transform 1 0 7312 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7646
timestamp 1018054153
transform 1 0 7328 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7648
timestamp 1018054153
transform 1 0 7344 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7650
timestamp 1018054153
transform 1 0 7360 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7652
timestamp 1018054153
transform 1 0 7376 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7654
timestamp 1018054153
transform 1 0 7392 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7656
timestamp 1018054153
transform 1 0 7408 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7658
timestamp 1018054153
transform 1 0 7424 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7660
timestamp 1018054153
transform 1 0 7440 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7662
timestamp 1018054153
transform 1 0 7456 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7664
timestamp 1018054153
transform 1 0 7472 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7666
timestamp 1018054153
transform 1 0 7488 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7668
timestamp 1018054153
transform 1 0 7504 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7670
timestamp 1018054153
transform 1 0 7520 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7672
timestamp 1018054153
transform 1 0 7536 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7674
timestamp 1018054153
transform 1 0 7552 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7676
timestamp 1018054153
transform 1 0 7568 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7678
timestamp 1018054153
transform 1 0 7584 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7680
timestamp 1018054153
transform 1 0 7600 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7682
timestamp 1018054153
transform 1 0 7616 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7684
timestamp 1018054153
transform 1 0 7632 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7686
timestamp 1018054153
transform 1 0 7648 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7688
timestamp 1018054153
transform 1 0 7664 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7690
timestamp 1018054153
transform 1 0 7680 0 -1 2880
box -16 -6 32 210
use FILL  FILL_7692
timestamp 1018054153
transform 1 0 7696 0 -1 2880
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_47
timestamp 1542725905
transform 1 0 7788 0 1 2680
box -48 -6 48 6
use FILL  FILL_7694
timestamp 1018054153
transform 1 0 7712 0 -1 2880
box -16 -6 32 210
use PADOUT  PADOUT_4
timestamp 1084294529
transform 0 1 8000 -1 0 3200
box -12 -6 606 2000
use M3_M2  M3_M2_126
timestamp 1542725905
transform 1 0 7848 0 1 2510
box -6 -6 6 6
use M3_M2  M3_M2_127
timestamp 1542725905
transform 1 0 8002 0 1 2510
box -6 -6 6 6
use mult_pad_VIA1  mult_pad_VIA1_48
timestamp 1542725905
transform 1 0 2092 0 1 2480
box -48 -6 48 6
use FILL  FILL_7695
timestamp 1018054153
transform 1 0 2272 0 1 2480
box -16 -6 32 210
use FILL  FILL_7697
timestamp 1018054153
transform 1 0 2288 0 1 2480
box -16 -6 32 210
use FILL  FILL_7699
timestamp 1018054153
transform 1 0 2304 0 1 2480
box -16 -6 32 210
use FILL  FILL_7701
timestamp 1018054153
transform 1 0 2320 0 1 2480
box -16 -6 32 210
use FILL  FILL_7703
timestamp 1018054153
transform 1 0 2336 0 1 2480
box -16 -6 32 210
use FILL  FILL_7705
timestamp 1018054153
transform 1 0 2352 0 1 2480
box -16 -6 32 210
use FILL  FILL_7707
timestamp 1018054153
transform 1 0 2368 0 1 2480
box -16 -6 32 210
use FILL  FILL_7709
timestamp 1018054153
transform 1 0 2384 0 1 2480
box -16 -6 32 210
use FILL  FILL_7711
timestamp 1018054153
transform 1 0 2400 0 1 2480
box -16 -6 32 210
use FILL  FILL_7713
timestamp 1018054153
transform 1 0 2416 0 1 2480
box -16 -6 32 210
use FILL  FILL_7715
timestamp 1018054153
transform 1 0 2432 0 1 2480
box -16 -6 32 210
use FILL  FILL_7717
timestamp 1018054153
transform 1 0 2448 0 1 2480
box -16 -6 32 210
use FILL  FILL_7719
timestamp 1018054153
transform 1 0 2464 0 1 2480
box -16 -6 32 210
use FILL  FILL_7721
timestamp 1018054153
transform 1 0 2480 0 1 2480
box -16 -6 32 210
use FILL  FILL_7723
timestamp 1018054153
transform 1 0 2496 0 1 2480
box -16 -6 32 210
use FILL  FILL_7725
timestamp 1018054153
transform 1 0 2512 0 1 2480
box -16 -6 32 210
use FILL  FILL_7727
timestamp 1018054153
transform 1 0 2528 0 1 2480
box -16 -6 32 210
use FILL  FILL_7729
timestamp 1018054153
transform 1 0 2544 0 1 2480
box -16 -6 32 210
use FILL  FILL_7731
timestamp 1018054153
transform 1 0 2560 0 1 2480
box -16 -6 32 210
use FILL  FILL_7733
timestamp 1018054153
transform 1 0 2576 0 1 2480
box -16 -6 32 210
use FILL  FILL_7735
timestamp 1018054153
transform 1 0 2592 0 1 2480
box -16 -6 32 210
use FILL  FILL_7737
timestamp 1018054153
transform 1 0 2608 0 1 2480
box -16 -6 32 210
use FILL  FILL_7739
timestamp 1018054153
transform 1 0 2624 0 1 2480
box -16 -6 32 210
use FILL  FILL_7741
timestamp 1018054153
transform 1 0 2640 0 1 2480
box -16 -6 32 210
use FILL  FILL_7743
timestamp 1018054153
transform 1 0 2656 0 1 2480
box -16 -6 32 210
use FILL  FILL_7745
timestamp 1018054153
transform 1 0 2672 0 1 2480
box -16 -6 32 210
use FILL  FILL_7747
timestamp 1018054153
transform 1 0 2688 0 1 2480
box -16 -6 32 210
use FILL  FILL_7749
timestamp 1018054153
transform 1 0 2704 0 1 2480
box -16 -6 32 210
use FILL  FILL_7751
timestamp 1018054153
transform 1 0 2720 0 1 2480
box -16 -6 32 210
use FILL  FILL_7753
timestamp 1018054153
transform 1 0 2736 0 1 2480
box -16 -6 32 210
use FILL  FILL_7755
timestamp 1018054153
transform 1 0 2752 0 1 2480
box -16 -6 32 210
use FILL  FILL_7757
timestamp 1018054153
transform 1 0 2768 0 1 2480
box -16 -6 32 210
use FILL  FILL_7759
timestamp 1018054153
transform 1 0 2784 0 1 2480
box -16 -6 32 210
use FILL  FILL_7761
timestamp 1018054153
transform 1 0 2800 0 1 2480
box -16 -6 32 210
use FILL  FILL_7763
timestamp 1018054153
transform 1 0 2816 0 1 2480
box -16 -6 32 210
use FILL  FILL_7765
timestamp 1018054153
transform 1 0 2832 0 1 2480
box -16 -6 32 210
use FILL  FILL_7767
timestamp 1018054153
transform 1 0 2848 0 1 2480
box -16 -6 32 210
use FILL  FILL_7769
timestamp 1018054153
transform 1 0 2864 0 1 2480
box -16 -6 32 210
use FILL  FILL_7771
timestamp 1018054153
transform 1 0 2880 0 1 2480
box -16 -6 32 210
use FILL  FILL_7773
timestamp 1018054153
transform 1 0 2896 0 1 2480
box -16 -6 32 210
use FILL  FILL_7775
timestamp 1018054153
transform 1 0 2912 0 1 2480
box -16 -6 32 210
use FILL  FILL_7777
timestamp 1018054153
transform 1 0 2928 0 1 2480
box -16 -6 32 210
use FILL  FILL_7779
timestamp 1018054153
transform 1 0 2944 0 1 2480
box -16 -6 32 210
use FILL  FILL_7781
timestamp 1018054153
transform 1 0 2960 0 1 2480
box -16 -6 32 210
use FILL  FILL_7783
timestamp 1018054153
transform 1 0 2976 0 1 2480
box -16 -6 32 210
use FILL  FILL_7785
timestamp 1018054153
transform 1 0 2992 0 1 2480
box -16 -6 32 210
use FILL  FILL_7787
timestamp 1018054153
transform 1 0 3008 0 1 2480
box -16 -6 32 210
use FILL  FILL_7789
timestamp 1018054153
transform 1 0 3024 0 1 2480
box -16 -6 32 210
use FILL  FILL_7791
timestamp 1018054153
transform 1 0 3040 0 1 2480
box -16 -6 32 210
use FILL  FILL_7793
timestamp 1018054153
transform 1 0 3056 0 1 2480
box -16 -6 32 210
use FILL  FILL_7795
timestamp 1018054153
transform 1 0 3072 0 1 2480
box -16 -6 32 210
use FILL  FILL_7797
timestamp 1018054153
transform 1 0 3088 0 1 2480
box -16 -6 32 210
use FILL  FILL_7799
timestamp 1018054153
transform 1 0 3104 0 1 2480
box -16 -6 32 210
use FILL  FILL_7801
timestamp 1018054153
transform 1 0 3120 0 1 2480
box -16 -6 32 210
use FILL  FILL_7803
timestamp 1018054153
transform 1 0 3136 0 1 2480
box -16 -6 32 210
use FILL  FILL_7805
timestamp 1018054153
transform 1 0 3152 0 1 2480
box -16 -6 32 210
use FILL  FILL_7807
timestamp 1018054153
transform 1 0 3168 0 1 2480
box -16 -6 32 210
use FILL  FILL_7809
timestamp 1018054153
transform 1 0 3184 0 1 2480
box -16 -6 32 210
use FILL  FILL_7811
timestamp 1018054153
transform 1 0 3200 0 1 2480
box -16 -6 32 210
use FILL  FILL_7813
timestamp 1018054153
transform 1 0 3216 0 1 2480
box -16 -6 32 210
use FILL  FILL_7815
timestamp 1018054153
transform 1 0 3232 0 1 2480
box -16 -6 32 210
use FILL  FILL_7817
timestamp 1018054153
transform 1 0 3248 0 1 2480
box -16 -6 32 210
use FILL  FILL_7819
timestamp 1018054153
transform 1 0 3264 0 1 2480
box -16 -6 32 210
use FILL  FILL_7821
timestamp 1018054153
transform 1 0 3280 0 1 2480
box -16 -6 32 210
use FILL  FILL_7823
timestamp 1018054153
transform 1 0 3296 0 1 2480
box -16 -6 32 210
use FILL  FILL_7825
timestamp 1018054153
transform 1 0 3312 0 1 2480
box -16 -6 32 210
use FILL  FILL_7827
timestamp 1018054153
transform 1 0 3328 0 1 2480
box -16 -6 32 210
use FILL  FILL_7829
timestamp 1018054153
transform 1 0 3344 0 1 2480
box -16 -6 32 210
use FILL  FILL_7831
timestamp 1018054153
transform 1 0 3360 0 1 2480
box -16 -6 32 210
use FILL  FILL_7833
timestamp 1018054153
transform 1 0 3376 0 1 2480
box -16 -6 32 210
use FILL  FILL_7835
timestamp 1018054153
transform 1 0 3392 0 1 2480
box -16 -6 32 210
use FILL  FILL_7837
timestamp 1018054153
transform 1 0 3408 0 1 2480
box -16 -6 32 210
use FILL  FILL_7839
timestamp 1018054153
transform 1 0 3424 0 1 2480
box -16 -6 32 210
use FILL  FILL_7841
timestamp 1018054153
transform 1 0 3440 0 1 2480
box -16 -6 32 210
use FILL  FILL_7843
timestamp 1018054153
transform 1 0 3456 0 1 2480
box -16 -6 32 210
use FILL  FILL_7845
timestamp 1018054153
transform 1 0 3472 0 1 2480
box -16 -6 32 210
use FILL  FILL_7847
timestamp 1018054153
transform 1 0 3488 0 1 2480
box -16 -6 32 210
use FILL  FILL_7849
timestamp 1018054153
transform 1 0 3504 0 1 2480
box -16 -6 32 210
use FILL  FILL_7851
timestamp 1018054153
transform 1 0 3520 0 1 2480
box -16 -6 32 210
use FILL  FILL_7853
timestamp 1018054153
transform 1 0 3536 0 1 2480
box -16 -6 32 210
use FILL  FILL_7855
timestamp 1018054153
transform 1 0 3552 0 1 2480
box -16 -6 32 210
use FILL  FILL_7857
timestamp 1018054153
transform 1 0 3568 0 1 2480
box -16 -6 32 210
use FILL  FILL_7859
timestamp 1018054153
transform 1 0 3584 0 1 2480
box -16 -6 32 210
use FILL  FILL_7861
timestamp 1018054153
transform 1 0 3600 0 1 2480
box -16 -6 32 210
use FILL  FILL_7863
timestamp 1018054153
transform 1 0 3616 0 1 2480
box -16 -6 32 210
use FILL  FILL_7865
timestamp 1018054153
transform 1 0 3632 0 1 2480
box -16 -6 32 210
use FILL  FILL_7867
timestamp 1018054153
transform 1 0 3648 0 1 2480
box -16 -6 32 210
use FILL  FILL_7869
timestamp 1018054153
transform 1 0 3664 0 1 2480
box -16 -6 32 210
use FILL  FILL_7871
timestamp 1018054153
transform 1 0 3680 0 1 2480
box -16 -6 32 210
use FILL  FILL_7873
timestamp 1018054153
transform 1 0 3696 0 1 2480
box -16 -6 32 210
use FILL  FILL_7875
timestamp 1018054153
transform 1 0 3712 0 1 2480
box -16 -6 32 210
use FILL  FILL_7877
timestamp 1018054153
transform 1 0 3728 0 1 2480
box -16 -6 32 210
use FILL  FILL_7879
timestamp 1018054153
transform 1 0 3744 0 1 2480
box -16 -6 32 210
use FILL  FILL_7881
timestamp 1018054153
transform 1 0 3760 0 1 2480
box -16 -6 32 210
use FILL  FILL_7883
timestamp 1018054153
transform 1 0 3776 0 1 2480
box -16 -6 32 210
use FILL  FILL_7885
timestamp 1018054153
transform 1 0 3792 0 1 2480
box -16 -6 32 210
use FILL  FILL_7887
timestamp 1018054153
transform 1 0 3808 0 1 2480
box -16 -6 32 210
use FILL  FILL_7889
timestamp 1018054153
transform 1 0 3824 0 1 2480
box -16 -6 32 210
use FILL  FILL_7891
timestamp 1018054153
transform 1 0 3840 0 1 2480
box -16 -6 32 210
use FILL  FILL_7893
timestamp 1018054153
transform 1 0 3856 0 1 2480
box -16 -6 32 210
use FILL  FILL_7895
timestamp 1018054153
transform 1 0 3872 0 1 2480
box -16 -6 32 210
use FILL  FILL_7897
timestamp 1018054153
transform 1 0 3888 0 1 2480
box -16 -6 32 210
use FILL  FILL_7899
timestamp 1018054153
transform 1 0 3904 0 1 2480
box -16 -6 32 210
use FILL  FILL_7901
timestamp 1018054153
transform 1 0 3920 0 1 2480
box -16 -6 32 210
use FILL  FILL_7903
timestamp 1018054153
transform 1 0 3936 0 1 2480
box -16 -6 32 210
use FILL  FILL_7905
timestamp 1018054153
transform 1 0 3952 0 1 2480
box -16 -6 32 210
use FILL  FILL_7907
timestamp 1018054153
transform 1 0 3968 0 1 2480
box -16 -6 32 210
use FILL  FILL_7909
timestamp 1018054153
transform 1 0 3984 0 1 2480
box -16 -6 32 210
use FILL  FILL_7911
timestamp 1018054153
transform 1 0 4000 0 1 2480
box -16 -6 32 210
use FILL  FILL_7913
timestamp 1018054153
transform 1 0 4016 0 1 2480
box -16 -6 32 210
use FILL  FILL_7915
timestamp 1018054153
transform 1 0 4032 0 1 2480
box -16 -6 32 210
use FILL  FILL_7917
timestamp 1018054153
transform 1 0 4048 0 1 2480
box -16 -6 32 210
use FILL  FILL_7919
timestamp 1018054153
transform 1 0 4064 0 1 2480
box -16 -6 32 210
use FILL  FILL_7921
timestamp 1018054153
transform 1 0 4080 0 1 2480
box -16 -6 32 210
use FILL  FILL_7923
timestamp 1018054153
transform 1 0 4096 0 1 2480
box -16 -6 32 210
use FILL  FILL_7925
timestamp 1018054153
transform 1 0 4112 0 1 2480
box -16 -6 32 210
use FILL  FILL_7927
timestamp 1018054153
transform 1 0 4128 0 1 2480
box -16 -6 32 210
use FILL  FILL_7929
timestamp 1018054153
transform 1 0 4144 0 1 2480
box -16 -6 32 210
use FILL  FILL_7931
timestamp 1018054153
transform 1 0 4160 0 1 2480
box -16 -6 32 210
use FILL  FILL_7933
timestamp 1018054153
transform 1 0 4176 0 1 2480
box -16 -6 32 210
use FILL  FILL_7935
timestamp 1018054153
transform 1 0 4192 0 1 2480
box -16 -6 32 210
use FILL  FILL_7937
timestamp 1018054153
transform 1 0 4208 0 1 2480
box -16 -6 32 210
use FILL  FILL_7939
timestamp 1018054153
transform 1 0 4224 0 1 2480
box -16 -6 32 210
use FILL  FILL_7941
timestamp 1018054153
transform 1 0 4240 0 1 2480
box -16 -6 32 210
use FILL  FILL_7943
timestamp 1018054153
transform 1 0 4256 0 1 2480
box -16 -6 32 210
use FILL  FILL_7945
timestamp 1018054153
transform 1 0 4272 0 1 2480
box -16 -6 32 210
use FILL  FILL_7947
timestamp 1018054153
transform 1 0 4288 0 1 2480
box -16 -6 32 210
use FILL  FILL_7949
timestamp 1018054153
transform 1 0 4304 0 1 2480
box -16 -6 32 210
use FILL  FILL_7951
timestamp 1018054153
transform 1 0 4320 0 1 2480
box -16 -6 32 210
use FILL  FILL_7953
timestamp 1018054153
transform 1 0 4336 0 1 2480
box -16 -6 32 210
use FILL  FILL_7955
timestamp 1018054153
transform 1 0 4352 0 1 2480
box -16 -6 32 210
use FILL  FILL_7957
timestamp 1018054153
transform 1 0 4368 0 1 2480
box -16 -6 32 210
use FILL  FILL_7959
timestamp 1018054153
transform 1 0 4384 0 1 2480
box -16 -6 32 210
use FILL  FILL_7961
timestamp 1018054153
transform 1 0 4400 0 1 2480
box -16 -6 32 210
use FILL  FILL_7963
timestamp 1018054153
transform 1 0 4416 0 1 2480
box -16 -6 32 210
use FILL  FILL_7965
timestamp 1018054153
transform 1 0 4432 0 1 2480
box -16 -6 32 210
use FILL  FILL_7967
timestamp 1018054153
transform 1 0 4448 0 1 2480
box -16 -6 32 210
use FILL  FILL_7969
timestamp 1018054153
transform 1 0 4464 0 1 2480
box -16 -6 32 210
use FILL  FILL_7971
timestamp 1018054153
transform 1 0 4480 0 1 2480
box -16 -6 32 210
use FILL  FILL_7973
timestamp 1018054153
transform 1 0 4496 0 1 2480
box -16 -6 32 210
use FILL  FILL_7975
timestamp 1018054153
transform 1 0 4512 0 1 2480
box -16 -6 32 210
use FILL  FILL_7977
timestamp 1018054153
transform 1 0 4528 0 1 2480
box -16 -6 32 210
use FILL  FILL_7979
timestamp 1018054153
transform 1 0 4544 0 1 2480
box -16 -6 32 210
use FILL  FILL_7981
timestamp 1018054153
transform 1 0 4560 0 1 2480
box -16 -6 32 210
use FILL  FILL_7983
timestamp 1018054153
transform 1 0 4576 0 1 2480
box -16 -6 32 210
use FILL  FILL_7985
timestamp 1018054153
transform 1 0 4592 0 1 2480
box -16 -6 32 210
use FILL  FILL_7987
timestamp 1018054153
transform 1 0 4608 0 1 2480
box -16 -6 32 210
use FILL  FILL_7989
timestamp 1018054153
transform 1 0 4624 0 1 2480
box -16 -6 32 210
use FILL  FILL_7991
timestamp 1018054153
transform 1 0 4640 0 1 2480
box -16 -6 32 210
use FILL  FILL_7993
timestamp 1018054153
transform 1 0 4656 0 1 2480
box -16 -6 32 210
use FILL  FILL_7995
timestamp 1018054153
transform 1 0 4672 0 1 2480
box -16 -6 32 210
use FILL  FILL_7997
timestamp 1018054153
transform 1 0 4688 0 1 2480
box -16 -6 32 210
use FILL  FILL_7999
timestamp 1018054153
transform 1 0 4704 0 1 2480
box -16 -6 32 210
use FILL  FILL_8001
timestamp 1018054153
transform 1 0 4720 0 1 2480
box -16 -6 32 210
use FILL  FILL_8003
timestamp 1018054153
transform 1 0 4736 0 1 2480
box -16 -6 32 210
use FILL  FILL_8005
timestamp 1018054153
transform 1 0 4752 0 1 2480
box -16 -6 32 210
use FILL  FILL_8007
timestamp 1018054153
transform 1 0 4768 0 1 2480
box -16 -6 32 210
use FILL  FILL_8009
timestamp 1018054153
transform 1 0 4784 0 1 2480
box -16 -6 32 210
use FILL  FILL_8011
timestamp 1018054153
transform 1 0 4800 0 1 2480
box -16 -6 32 210
use FILL  FILL_8013
timestamp 1018054153
transform 1 0 4816 0 1 2480
box -16 -6 32 210
use FILL  FILL_8015
timestamp 1018054153
transform 1 0 4832 0 1 2480
box -16 -6 32 210
use FILL  FILL_8017
timestamp 1018054153
transform 1 0 4848 0 1 2480
box -16 -6 32 210
use FILL  FILL_8019
timestamp 1018054153
transform 1 0 4864 0 1 2480
box -16 -6 32 210
use FILL  FILL_8021
timestamp 1018054153
transform 1 0 4880 0 1 2480
box -16 -6 32 210
use FILL  FILL_8023
timestamp 1018054153
transform 1 0 4896 0 1 2480
box -16 -6 32 210
use FILL  FILL_8025
timestamp 1018054153
transform 1 0 4912 0 1 2480
box -16 -6 32 210
use FILL  FILL_8027
timestamp 1018054153
transform 1 0 4928 0 1 2480
box -16 -6 32 210
use FILL  FILL_8029
timestamp 1018054153
transform 1 0 4944 0 1 2480
box -16 -6 32 210
use FILL  FILL_8031
timestamp 1018054153
transform 1 0 4960 0 1 2480
box -16 -6 32 210
use FILL  FILL_8033
timestamp 1018054153
transform 1 0 4976 0 1 2480
box -16 -6 32 210
use FILL  FILL_8035
timestamp 1018054153
transform 1 0 4992 0 1 2480
box -16 -6 32 210
use FILL  FILL_8037
timestamp 1018054153
transform 1 0 5008 0 1 2480
box -16 -6 32 210
use FILL  FILL_8039
timestamp 1018054153
transform 1 0 5024 0 1 2480
box -16 -6 32 210
use FILL  FILL_8041
timestamp 1018054153
transform 1 0 5040 0 1 2480
box -16 -6 32 210
use FILL  FILL_8043
timestamp 1018054153
transform 1 0 5056 0 1 2480
box -16 -6 32 210
use FILL  FILL_8045
timestamp 1018054153
transform 1 0 5072 0 1 2480
box -16 -6 32 210
use FILL  FILL_8047
timestamp 1018054153
transform 1 0 5088 0 1 2480
box -16 -6 32 210
use FILL  FILL_8049
timestamp 1018054153
transform 1 0 5104 0 1 2480
box -16 -6 32 210
use FILL  FILL_8051
timestamp 1018054153
transform 1 0 5120 0 1 2480
box -16 -6 32 210
use FILL  FILL_8053
timestamp 1018054153
transform 1 0 5136 0 1 2480
box -16 -6 32 210
use FILL  FILL_8055
timestamp 1018054153
transform 1 0 5152 0 1 2480
box -16 -6 32 210
use FILL  FILL_8057
timestamp 1018054153
transform 1 0 5168 0 1 2480
box -16 -6 32 210
use FILL  FILL_8059
timestamp 1018054153
transform 1 0 5184 0 1 2480
box -16 -6 32 210
use FILL  FILL_8061
timestamp 1018054153
transform 1 0 5200 0 1 2480
box -16 -6 32 210
use FILL  FILL_8063
timestamp 1018054153
transform 1 0 5216 0 1 2480
box -16 -6 32 210
use FILL  FILL_8065
timestamp 1018054153
transform 1 0 5232 0 1 2480
box -16 -6 32 210
use FILL  FILL_8067
timestamp 1018054153
transform 1 0 5248 0 1 2480
box -16 -6 32 210
use FILL  FILL_8069
timestamp 1018054153
transform 1 0 5264 0 1 2480
box -16 -6 32 210
use FILL  FILL_8071
timestamp 1018054153
transform 1 0 5280 0 1 2480
box -16 -6 32 210
use FILL  FILL_8073
timestamp 1018054153
transform 1 0 5296 0 1 2480
box -16 -6 32 210
use FILL  FILL_8075
timestamp 1018054153
transform 1 0 5312 0 1 2480
box -16 -6 32 210
use FILL  FILL_8077
timestamp 1018054153
transform 1 0 5328 0 1 2480
box -16 -6 32 210
use FILL  FILL_8079
timestamp 1018054153
transform 1 0 5344 0 1 2480
box -16 -6 32 210
use FILL  FILL_8081
timestamp 1018054153
transform 1 0 5360 0 1 2480
box -16 -6 32 210
use FILL  FILL_8083
timestamp 1018054153
transform 1 0 5376 0 1 2480
box -16 -6 32 210
use FILL  FILL_8085
timestamp 1018054153
transform 1 0 5392 0 1 2480
box -16 -6 32 210
use FILL  FILL_8087
timestamp 1018054153
transform 1 0 5408 0 1 2480
box -16 -6 32 210
use FILL  FILL_8089
timestamp 1018054153
transform 1 0 5424 0 1 2480
box -16 -6 32 210
use FILL  FILL_8091
timestamp 1018054153
transform 1 0 5440 0 1 2480
box -16 -6 32 210
use FILL  FILL_8093
timestamp 1018054153
transform 1 0 5456 0 1 2480
box -16 -6 32 210
use FILL  FILL_8095
timestamp 1018054153
transform 1 0 5472 0 1 2480
box -16 -6 32 210
use FILL  FILL_8097
timestamp 1018054153
transform 1 0 5488 0 1 2480
box -16 -6 32 210
use FILL  FILL_8099
timestamp 1018054153
transform 1 0 5504 0 1 2480
box -16 -6 32 210
use FILL  FILL_8101
timestamp 1018054153
transform 1 0 5520 0 1 2480
box -16 -6 32 210
use FILL  FILL_8103
timestamp 1018054153
transform 1 0 5536 0 1 2480
box -16 -6 32 210
use FILL  FILL_8105
timestamp 1018054153
transform 1 0 5552 0 1 2480
box -16 -6 32 210
use FILL  FILL_8107
timestamp 1018054153
transform 1 0 5568 0 1 2480
box -16 -6 32 210
use FILL  FILL_8109
timestamp 1018054153
transform 1 0 5584 0 1 2480
box -16 -6 32 210
use FILL  FILL_8111
timestamp 1018054153
transform 1 0 5600 0 1 2480
box -16 -6 32 210
use FILL  FILL_8113
timestamp 1018054153
transform 1 0 5616 0 1 2480
box -16 -6 32 210
use FILL  FILL_8115
timestamp 1018054153
transform 1 0 5632 0 1 2480
box -16 -6 32 210
use FILL  FILL_8117
timestamp 1018054153
transform 1 0 5648 0 1 2480
box -16 -6 32 210
use FILL  FILL_8119
timestamp 1018054153
transform 1 0 5664 0 1 2480
box -16 -6 32 210
use FILL  FILL_8121
timestamp 1018054153
transform 1 0 5680 0 1 2480
box -16 -6 32 210
use FILL  FILL_8123
timestamp 1018054153
transform 1 0 5696 0 1 2480
box -16 -6 32 210
use FILL  FILL_8125
timestamp 1018054153
transform 1 0 5712 0 1 2480
box -16 -6 32 210
use FILL  FILL_8127
timestamp 1018054153
transform 1 0 5728 0 1 2480
box -16 -6 32 210
use FILL  FILL_8129
timestamp 1018054153
transform 1 0 5744 0 1 2480
box -16 -6 32 210
use FILL  FILL_8131
timestamp 1018054153
transform 1 0 5760 0 1 2480
box -16 -6 32 210
use FILL  FILL_8133
timestamp 1018054153
transform 1 0 5776 0 1 2480
box -16 -6 32 210
use FILL  FILL_8135
timestamp 1018054153
transform 1 0 5792 0 1 2480
box -16 -6 32 210
use FILL  FILL_8137
timestamp 1018054153
transform 1 0 5808 0 1 2480
box -16 -6 32 210
use FILL  FILL_8139
timestamp 1018054153
transform 1 0 5824 0 1 2480
box -16 -6 32 210
use FILL  FILL_8141
timestamp 1018054153
transform 1 0 5840 0 1 2480
box -16 -6 32 210
use FILL  FILL_8143
timestamp 1018054153
transform 1 0 5856 0 1 2480
box -16 -6 32 210
use FILL  FILL_8145
timestamp 1018054153
transform 1 0 5872 0 1 2480
box -16 -6 32 210
use FILL  FILL_8147
timestamp 1018054153
transform 1 0 5888 0 1 2480
box -16 -6 32 210
use FILL  FILL_8149
timestamp 1018054153
transform 1 0 5904 0 1 2480
box -16 -6 32 210
use FILL  FILL_8151
timestamp 1018054153
transform 1 0 5920 0 1 2480
box -16 -6 32 210
use FILL  FILL_8153
timestamp 1018054153
transform 1 0 5936 0 1 2480
box -16 -6 32 210
use FILL  FILL_8155
timestamp 1018054153
transform 1 0 5952 0 1 2480
box -16 -6 32 210
use FILL  FILL_8157
timestamp 1018054153
transform 1 0 5968 0 1 2480
box -16 -6 32 210
use FILL  FILL_8159
timestamp 1018054153
transform 1 0 5984 0 1 2480
box -16 -6 32 210
use FILL  FILL_8161
timestamp 1018054153
transform 1 0 6000 0 1 2480
box -16 -6 32 210
use FILL  FILL_8163
timestamp 1018054153
transform 1 0 6016 0 1 2480
box -16 -6 32 210
use FILL  FILL_8165
timestamp 1018054153
transform 1 0 6032 0 1 2480
box -16 -6 32 210
use FILL  FILL_8167
timestamp 1018054153
transform 1 0 6048 0 1 2480
box -16 -6 32 210
use FILL  FILL_8169
timestamp 1018054153
transform 1 0 6064 0 1 2480
box -16 -6 32 210
use FILL  FILL_8171
timestamp 1018054153
transform 1 0 6080 0 1 2480
box -16 -6 32 210
use FILL  FILL_8173
timestamp 1018054153
transform 1 0 6096 0 1 2480
box -16 -6 32 210
use FILL  FILL_8175
timestamp 1018054153
transform 1 0 6112 0 1 2480
box -16 -6 32 210
use FILL  FILL_8177
timestamp 1018054153
transform 1 0 6128 0 1 2480
box -16 -6 32 210
use FILL  FILL_8179
timestamp 1018054153
transform 1 0 6144 0 1 2480
box -16 -6 32 210
use FILL  FILL_8181
timestamp 1018054153
transform 1 0 6160 0 1 2480
box -16 -6 32 210
use FILL  FILL_8183
timestamp 1018054153
transform 1 0 6176 0 1 2480
box -16 -6 32 210
use FILL  FILL_8185
timestamp 1018054153
transform 1 0 6192 0 1 2480
box -16 -6 32 210
use FILL  FILL_8187
timestamp 1018054153
transform 1 0 6208 0 1 2480
box -16 -6 32 210
use FILL  FILL_8189
timestamp 1018054153
transform 1 0 6224 0 1 2480
box -16 -6 32 210
use FILL  FILL_8191
timestamp 1018054153
transform 1 0 6240 0 1 2480
box -16 -6 32 210
use FILL  FILL_8193
timestamp 1018054153
transform 1 0 6256 0 1 2480
box -16 -6 32 210
use FILL  FILL_8195
timestamp 1018054153
transform 1 0 6272 0 1 2480
box -16 -6 32 210
use FILL  FILL_8197
timestamp 1018054153
transform 1 0 6288 0 1 2480
box -16 -6 32 210
use FILL  FILL_8199
timestamp 1018054153
transform 1 0 6304 0 1 2480
box -16 -6 32 210
use FILL  FILL_8201
timestamp 1018054153
transform 1 0 6320 0 1 2480
box -16 -6 32 210
use FILL  FILL_8203
timestamp 1018054153
transform 1 0 6336 0 1 2480
box -16 -6 32 210
use FILL  FILL_8205
timestamp 1018054153
transform 1 0 6352 0 1 2480
box -16 -6 32 210
use FILL  FILL_8207
timestamp 1018054153
transform 1 0 6368 0 1 2480
box -16 -6 32 210
use FILL  FILL_8209
timestamp 1018054153
transform 1 0 6384 0 1 2480
box -16 -6 32 210
use FILL  FILL_8211
timestamp 1018054153
transform 1 0 6400 0 1 2480
box -16 -6 32 210
use FILL  FILL_8213
timestamp 1018054153
transform 1 0 6416 0 1 2480
box -16 -6 32 210
use FILL  FILL_8215
timestamp 1018054153
transform 1 0 6432 0 1 2480
box -16 -6 32 210
use FILL  FILL_8217
timestamp 1018054153
transform 1 0 6448 0 1 2480
box -16 -6 32 210
use FILL  FILL_8219
timestamp 1018054153
transform 1 0 6464 0 1 2480
box -16 -6 32 210
use FILL  FILL_8221
timestamp 1018054153
transform 1 0 6480 0 1 2480
box -16 -6 32 210
use FILL  FILL_8223
timestamp 1018054153
transform 1 0 6496 0 1 2480
box -16 -6 32 210
use FILL  FILL_8225
timestamp 1018054153
transform 1 0 6512 0 1 2480
box -16 -6 32 210
use FILL  FILL_8227
timestamp 1018054153
transform 1 0 6528 0 1 2480
box -16 -6 32 210
use FILL  FILL_8229
timestamp 1018054153
transform 1 0 6544 0 1 2480
box -16 -6 32 210
use FILL  FILL_8231
timestamp 1018054153
transform 1 0 6560 0 1 2480
box -16 -6 32 210
use FILL  FILL_8233
timestamp 1018054153
transform 1 0 6576 0 1 2480
box -16 -6 32 210
use FILL  FILL_8235
timestamp 1018054153
transform 1 0 6592 0 1 2480
box -16 -6 32 210
use FILL  FILL_8237
timestamp 1018054153
transform 1 0 6608 0 1 2480
box -16 -6 32 210
use FILL  FILL_8239
timestamp 1018054153
transform 1 0 6624 0 1 2480
box -16 -6 32 210
use FILL  FILL_8241
timestamp 1018054153
transform 1 0 6640 0 1 2480
box -16 -6 32 210
use FILL  FILL_8243
timestamp 1018054153
transform 1 0 6656 0 1 2480
box -16 -6 32 210
use FILL  FILL_8245
timestamp 1018054153
transform 1 0 6672 0 1 2480
box -16 -6 32 210
use FILL  FILL_8247
timestamp 1018054153
transform 1 0 6688 0 1 2480
box -16 -6 32 210
use FILL  FILL_8249
timestamp 1018054153
transform 1 0 6704 0 1 2480
box -16 -6 32 210
use FILL  FILL_8251
timestamp 1018054153
transform 1 0 6720 0 1 2480
box -16 -6 32 210
use FILL  FILL_8253
timestamp 1018054153
transform 1 0 6736 0 1 2480
box -16 -6 32 210
use FILL  FILL_8255
timestamp 1018054153
transform 1 0 6752 0 1 2480
box -16 -6 32 210
use FILL  FILL_8257
timestamp 1018054153
transform 1 0 6768 0 1 2480
box -16 -6 32 210
use FILL  FILL_8259
timestamp 1018054153
transform 1 0 6784 0 1 2480
box -16 -6 32 210
use FILL  FILL_8261
timestamp 1018054153
transform 1 0 6800 0 1 2480
box -16 -6 32 210
use FILL  FILL_8263
timestamp 1018054153
transform 1 0 6816 0 1 2480
box -16 -6 32 210
use FILL  FILL_8265
timestamp 1018054153
transform 1 0 6832 0 1 2480
box -16 -6 32 210
use FILL  FILL_8267
timestamp 1018054153
transform 1 0 6848 0 1 2480
box -16 -6 32 210
use FILL  FILL_8269
timestamp 1018054153
transform 1 0 6864 0 1 2480
box -16 -6 32 210
use FILL  FILL_8271
timestamp 1018054153
transform 1 0 6880 0 1 2480
box -16 -6 32 210
use FILL  FILL_8273
timestamp 1018054153
transform 1 0 6896 0 1 2480
box -16 -6 32 210
use FILL  FILL_8275
timestamp 1018054153
transform 1 0 6912 0 1 2480
box -16 -6 32 210
use FILL  FILL_8277
timestamp 1018054153
transform 1 0 6928 0 1 2480
box -16 -6 32 210
use FILL  FILL_8279
timestamp 1018054153
transform 1 0 6944 0 1 2480
box -16 -6 32 210
use FILL  FILL_8281
timestamp 1018054153
transform 1 0 6960 0 1 2480
box -16 -6 32 210
use FILL  FILL_8283
timestamp 1018054153
transform 1 0 6976 0 1 2480
box -16 -6 32 210
use FILL  FILL_8285
timestamp 1018054153
transform 1 0 6992 0 1 2480
box -16 -6 32 210
use FILL  FILL_8287
timestamp 1018054153
transform 1 0 7008 0 1 2480
box -16 -6 32 210
use FILL  FILL_8289
timestamp 1018054153
transform 1 0 7024 0 1 2480
box -16 -6 32 210
use FILL  FILL_8291
timestamp 1018054153
transform 1 0 7040 0 1 2480
box -16 -6 32 210
use FILL  FILL_8293
timestamp 1018054153
transform 1 0 7056 0 1 2480
box -16 -6 32 210
use FILL  FILL_8295
timestamp 1018054153
transform 1 0 7072 0 1 2480
box -16 -6 32 210
use FILL  FILL_8297
timestamp 1018054153
transform 1 0 7088 0 1 2480
box -16 -6 32 210
use FILL  FILL_8299
timestamp 1018054153
transform 1 0 7104 0 1 2480
box -16 -6 32 210
use FILL  FILL_8301
timestamp 1018054153
transform 1 0 7120 0 1 2480
box -16 -6 32 210
use FILL  FILL_8303
timestamp 1018054153
transform 1 0 7136 0 1 2480
box -16 -6 32 210
use FILL  FILL_8305
timestamp 1018054153
transform 1 0 7152 0 1 2480
box -16 -6 32 210
use FILL  FILL_8307
timestamp 1018054153
transform 1 0 7168 0 1 2480
box -16 -6 32 210
use FILL  FILL_8309
timestamp 1018054153
transform 1 0 7184 0 1 2480
box -16 -6 32 210
use FILL  FILL_8311
timestamp 1018054153
transform 1 0 7200 0 1 2480
box -16 -6 32 210
use FILL  FILL_8313
timestamp 1018054153
transform 1 0 7216 0 1 2480
box -16 -6 32 210
use FILL  FILL_8315
timestamp 1018054153
transform 1 0 7232 0 1 2480
box -16 -6 32 210
use FILL  FILL_8317
timestamp 1018054153
transform 1 0 7248 0 1 2480
box -16 -6 32 210
use FILL  FILL_8319
timestamp 1018054153
transform 1 0 7264 0 1 2480
box -16 -6 32 210
use FILL  FILL_8321
timestamp 1018054153
transform 1 0 7280 0 1 2480
box -16 -6 32 210
use FILL  FILL_8323
timestamp 1018054153
transform 1 0 7296 0 1 2480
box -16 -6 32 210
use FILL  FILL_8325
timestamp 1018054153
transform 1 0 7312 0 1 2480
box -16 -6 32 210
use FILL  FILL_8327
timestamp 1018054153
transform 1 0 7328 0 1 2480
box -16 -6 32 210
use FILL  FILL_8329
timestamp 1018054153
transform 1 0 7344 0 1 2480
box -16 -6 32 210
use FILL  FILL_8331
timestamp 1018054153
transform 1 0 7360 0 1 2480
box -16 -6 32 210
use FILL  FILL_8333
timestamp 1018054153
transform 1 0 7376 0 1 2480
box -16 -6 32 210
use FILL  FILL_8335
timestamp 1018054153
transform 1 0 7392 0 1 2480
box -16 -6 32 210
use FILL  FILL_8337
timestamp 1018054153
transform 1 0 7408 0 1 2480
box -16 -6 32 210
use FILL  FILL_8339
timestamp 1018054153
transform 1 0 7424 0 1 2480
box -16 -6 32 210
use FILL  FILL_8341
timestamp 1018054153
transform 1 0 7440 0 1 2480
box -16 -6 32 210
use FILL  FILL_8343
timestamp 1018054153
transform 1 0 7456 0 1 2480
box -16 -6 32 210
use FILL  FILL_8345
timestamp 1018054153
transform 1 0 7472 0 1 2480
box -16 -6 32 210
use FILL  FILL_8347
timestamp 1018054153
transform 1 0 7488 0 1 2480
box -16 -6 32 210
use FILL  FILL_8349
timestamp 1018054153
transform 1 0 7504 0 1 2480
box -16 -6 32 210
use FILL  FILL_8351
timestamp 1018054153
transform 1 0 7520 0 1 2480
box -16 -6 32 210
use FILL  FILL_8353
timestamp 1018054153
transform 1 0 7536 0 1 2480
box -16 -6 32 210
use FILL  FILL_8355
timestamp 1018054153
transform 1 0 7552 0 1 2480
box -16 -6 32 210
use FILL  FILL_8357
timestamp 1018054153
transform 1 0 7568 0 1 2480
box -16 -6 32 210
use FILL  FILL_8359
timestamp 1018054153
transform 1 0 7584 0 1 2480
box -16 -6 32 210
use FILL  FILL_8361
timestamp 1018054153
transform 1 0 7600 0 1 2480
box -16 -6 32 210
use FILL  FILL_8363
timestamp 1018054153
transform 1 0 7616 0 1 2480
box -16 -6 32 210
use FILL  FILL_8365
timestamp 1018054153
transform 1 0 7632 0 1 2480
box -16 -6 32 210
use FILL  FILL_8367
timestamp 1018054153
transform 1 0 7648 0 1 2480
box -16 -6 32 210
use FILL  FILL_8369
timestamp 1018054153
transform 1 0 7664 0 1 2480
box -16 -6 32 210
use FILL  FILL_8371
timestamp 1018054153
transform 1 0 7680 0 1 2480
box -16 -6 32 210
use FILL  FILL_8373
timestamp 1018054153
transform 1 0 7696 0 1 2480
box -16 -6 32 210
use FILL  FILL_8375
timestamp 1018054153
transform 1 0 7712 0 1 2480
box -16 -6 32 210
use mult_pad_VIA1  mult_pad_VIA1_49
timestamp 1542725905
transform 1 0 7908 0 1 2480
box -48 -6 48 6
use mult_pad_VIA1  mult_pad_VIA1_50
timestamp 1542725905
transform 1 0 2212 0 1 2280
box -48 -6 48 6
use FILL  FILL_7696
timestamp 1018054153
transform 1 0 2272 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7698
timestamp 1018054153
transform 1 0 2288 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7700
timestamp 1018054153
transform 1 0 2304 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7702
timestamp 1018054153
transform 1 0 2320 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7704
timestamp 1018054153
transform 1 0 2336 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7706
timestamp 1018054153
transform 1 0 2352 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7708
timestamp 1018054153
transform 1 0 2368 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7710
timestamp 1018054153
transform 1 0 2384 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7712
timestamp 1018054153
transform 1 0 2400 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7714
timestamp 1018054153
transform 1 0 2416 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7716
timestamp 1018054153
transform 1 0 2432 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7718
timestamp 1018054153
transform 1 0 2448 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7720
timestamp 1018054153
transform 1 0 2464 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7722
timestamp 1018054153
transform 1 0 2480 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7724
timestamp 1018054153
transform 1 0 2496 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7726
timestamp 1018054153
transform 1 0 2512 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7728
timestamp 1018054153
transform 1 0 2528 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7730
timestamp 1018054153
transform 1 0 2544 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7732
timestamp 1018054153
transform 1 0 2560 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7734
timestamp 1018054153
transform 1 0 2576 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7736
timestamp 1018054153
transform 1 0 2592 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7738
timestamp 1018054153
transform 1 0 2608 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7740
timestamp 1018054153
transform 1 0 2624 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7742
timestamp 1018054153
transform 1 0 2640 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7744
timestamp 1018054153
transform 1 0 2656 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7746
timestamp 1018054153
transform 1 0 2672 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7748
timestamp 1018054153
transform 1 0 2688 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7750
timestamp 1018054153
transform 1 0 2704 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7752
timestamp 1018054153
transform 1 0 2720 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7754
timestamp 1018054153
transform 1 0 2736 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7756
timestamp 1018054153
transform 1 0 2752 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7758
timestamp 1018054153
transform 1 0 2768 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7760
timestamp 1018054153
transform 1 0 2784 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7762
timestamp 1018054153
transform 1 0 2800 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7764
timestamp 1018054153
transform 1 0 2816 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7766
timestamp 1018054153
transform 1 0 2832 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7768
timestamp 1018054153
transform 1 0 2848 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7770
timestamp 1018054153
transform 1 0 2864 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7772
timestamp 1018054153
transform 1 0 2880 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7774
timestamp 1018054153
transform 1 0 2896 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7776
timestamp 1018054153
transform 1 0 2912 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7778
timestamp 1018054153
transform 1 0 2928 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7780
timestamp 1018054153
transform 1 0 2944 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7782
timestamp 1018054153
transform 1 0 2960 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7784
timestamp 1018054153
transform 1 0 2976 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7786
timestamp 1018054153
transform 1 0 2992 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7788
timestamp 1018054153
transform 1 0 3008 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7790
timestamp 1018054153
transform 1 0 3024 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7792
timestamp 1018054153
transform 1 0 3040 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7794
timestamp 1018054153
transform 1 0 3056 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7796
timestamp 1018054153
transform 1 0 3072 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7798
timestamp 1018054153
transform 1 0 3088 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7800
timestamp 1018054153
transform 1 0 3104 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7802
timestamp 1018054153
transform 1 0 3120 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7804
timestamp 1018054153
transform 1 0 3136 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7806
timestamp 1018054153
transform 1 0 3152 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7808
timestamp 1018054153
transform 1 0 3168 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7810
timestamp 1018054153
transform 1 0 3184 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7812
timestamp 1018054153
transform 1 0 3200 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7814
timestamp 1018054153
transform 1 0 3216 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7816
timestamp 1018054153
transform 1 0 3232 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7818
timestamp 1018054153
transform 1 0 3248 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7820
timestamp 1018054153
transform 1 0 3264 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7822
timestamp 1018054153
transform 1 0 3280 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7824
timestamp 1018054153
transform 1 0 3296 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7826
timestamp 1018054153
transform 1 0 3312 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7828
timestamp 1018054153
transform 1 0 3328 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7830
timestamp 1018054153
transform 1 0 3344 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7832
timestamp 1018054153
transform 1 0 3360 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7834
timestamp 1018054153
transform 1 0 3376 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7836
timestamp 1018054153
transform 1 0 3392 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7838
timestamp 1018054153
transform 1 0 3408 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7840
timestamp 1018054153
transform 1 0 3424 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7842
timestamp 1018054153
transform 1 0 3440 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7844
timestamp 1018054153
transform 1 0 3456 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7846
timestamp 1018054153
transform 1 0 3472 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7848
timestamp 1018054153
transform 1 0 3488 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7850
timestamp 1018054153
transform 1 0 3504 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7852
timestamp 1018054153
transform 1 0 3520 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7854
timestamp 1018054153
transform 1 0 3536 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7856
timestamp 1018054153
transform 1 0 3552 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7858
timestamp 1018054153
transform 1 0 3568 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7860
timestamp 1018054153
transform 1 0 3584 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7862
timestamp 1018054153
transform 1 0 3600 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7864
timestamp 1018054153
transform 1 0 3616 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7866
timestamp 1018054153
transform 1 0 3632 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7868
timestamp 1018054153
transform 1 0 3648 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7870
timestamp 1018054153
transform 1 0 3664 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7872
timestamp 1018054153
transform 1 0 3680 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7874
timestamp 1018054153
transform 1 0 3696 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7876
timestamp 1018054153
transform 1 0 3712 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7878
timestamp 1018054153
transform 1 0 3728 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7880
timestamp 1018054153
transform 1 0 3744 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7882
timestamp 1018054153
transform 1 0 3760 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7884
timestamp 1018054153
transform 1 0 3776 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7886
timestamp 1018054153
transform 1 0 3792 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7888
timestamp 1018054153
transform 1 0 3808 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7890
timestamp 1018054153
transform 1 0 3824 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7892
timestamp 1018054153
transform 1 0 3840 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7894
timestamp 1018054153
transform 1 0 3856 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7896
timestamp 1018054153
transform 1 0 3872 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7898
timestamp 1018054153
transform 1 0 3888 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7900
timestamp 1018054153
transform 1 0 3904 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7902
timestamp 1018054153
transform 1 0 3920 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7904
timestamp 1018054153
transform 1 0 3936 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7906
timestamp 1018054153
transform 1 0 3952 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7908
timestamp 1018054153
transform 1 0 3968 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7910
timestamp 1018054153
transform 1 0 3984 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7912
timestamp 1018054153
transform 1 0 4000 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7914
timestamp 1018054153
transform 1 0 4016 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7916
timestamp 1018054153
transform 1 0 4032 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7918
timestamp 1018054153
transform 1 0 4048 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7920
timestamp 1018054153
transform 1 0 4064 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7922
timestamp 1018054153
transform 1 0 4080 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7924
timestamp 1018054153
transform 1 0 4096 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7926
timestamp 1018054153
transform 1 0 4112 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7928
timestamp 1018054153
transform 1 0 4128 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7930
timestamp 1018054153
transform 1 0 4144 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7932
timestamp 1018054153
transform 1 0 4160 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7934
timestamp 1018054153
transform 1 0 4176 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7936
timestamp 1018054153
transform 1 0 4192 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7938
timestamp 1018054153
transform 1 0 4208 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7940
timestamp 1018054153
transform 1 0 4224 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7942
timestamp 1018054153
transform 1 0 4240 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7944
timestamp 1018054153
transform 1 0 4256 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7946
timestamp 1018054153
transform 1 0 4272 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7948
timestamp 1018054153
transform 1 0 4288 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7950
timestamp 1018054153
transform 1 0 4304 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7952
timestamp 1018054153
transform 1 0 4320 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7954
timestamp 1018054153
transform 1 0 4336 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7956
timestamp 1018054153
transform 1 0 4352 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7958
timestamp 1018054153
transform 1 0 4368 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7960
timestamp 1018054153
transform 1 0 4384 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7962
timestamp 1018054153
transform 1 0 4400 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7964
timestamp 1018054153
transform 1 0 4416 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7966
timestamp 1018054153
transform 1 0 4432 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7968
timestamp 1018054153
transform 1 0 4448 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7970
timestamp 1018054153
transform 1 0 4464 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7972
timestamp 1018054153
transform 1 0 4480 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7974
timestamp 1018054153
transform 1 0 4496 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7976
timestamp 1018054153
transform 1 0 4512 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7978
timestamp 1018054153
transform 1 0 4528 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7980
timestamp 1018054153
transform 1 0 4544 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7982
timestamp 1018054153
transform 1 0 4560 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7984
timestamp 1018054153
transform 1 0 4576 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7986
timestamp 1018054153
transform 1 0 4592 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7988
timestamp 1018054153
transform 1 0 4608 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7990
timestamp 1018054153
transform 1 0 4624 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7992
timestamp 1018054153
transform 1 0 4640 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7994
timestamp 1018054153
transform 1 0 4656 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7996
timestamp 1018054153
transform 1 0 4672 0 -1 2480
box -16 -6 32 210
use FILL  FILL_7998
timestamp 1018054153
transform 1 0 4688 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8000
timestamp 1018054153
transform 1 0 4704 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8002
timestamp 1018054153
transform 1 0 4720 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8004
timestamp 1018054153
transform 1 0 4736 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8006
timestamp 1018054153
transform 1 0 4752 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8008
timestamp 1018054153
transform 1 0 4768 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8010
timestamp 1018054153
transform 1 0 4784 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8012
timestamp 1018054153
transform 1 0 4800 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8014
timestamp 1018054153
transform 1 0 4816 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8016
timestamp 1018054153
transform 1 0 4832 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8018
timestamp 1018054153
transform 1 0 4848 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8020
timestamp 1018054153
transform 1 0 4864 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8022
timestamp 1018054153
transform 1 0 4880 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8024
timestamp 1018054153
transform 1 0 4896 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8026
timestamp 1018054153
transform 1 0 4912 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8028
timestamp 1018054153
transform 1 0 4928 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8030
timestamp 1018054153
transform 1 0 4944 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8032
timestamp 1018054153
transform 1 0 4960 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8034
timestamp 1018054153
transform 1 0 4976 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8036
timestamp 1018054153
transform 1 0 4992 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8038
timestamp 1018054153
transform 1 0 5008 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8040
timestamp 1018054153
transform 1 0 5024 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8042
timestamp 1018054153
transform 1 0 5040 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8044
timestamp 1018054153
transform 1 0 5056 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8046
timestamp 1018054153
transform 1 0 5072 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8048
timestamp 1018054153
transform 1 0 5088 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8050
timestamp 1018054153
transform 1 0 5104 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8052
timestamp 1018054153
transform 1 0 5120 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8054
timestamp 1018054153
transform 1 0 5136 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8056
timestamp 1018054153
transform 1 0 5152 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8058
timestamp 1018054153
transform 1 0 5168 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8060
timestamp 1018054153
transform 1 0 5184 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8062
timestamp 1018054153
transform 1 0 5200 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8064
timestamp 1018054153
transform 1 0 5216 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8066
timestamp 1018054153
transform 1 0 5232 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8068
timestamp 1018054153
transform 1 0 5248 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8070
timestamp 1018054153
transform 1 0 5264 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8072
timestamp 1018054153
transform 1 0 5280 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8074
timestamp 1018054153
transform 1 0 5296 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8076
timestamp 1018054153
transform 1 0 5312 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8078
timestamp 1018054153
transform 1 0 5328 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8080
timestamp 1018054153
transform 1 0 5344 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8082
timestamp 1018054153
transform 1 0 5360 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8084
timestamp 1018054153
transform 1 0 5376 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8086
timestamp 1018054153
transform 1 0 5392 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8088
timestamp 1018054153
transform 1 0 5408 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8090
timestamp 1018054153
transform 1 0 5424 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8092
timestamp 1018054153
transform 1 0 5440 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8094
timestamp 1018054153
transform 1 0 5456 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8096
timestamp 1018054153
transform 1 0 5472 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8098
timestamp 1018054153
transform 1 0 5488 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8100
timestamp 1018054153
transform 1 0 5504 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8102
timestamp 1018054153
transform 1 0 5520 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8104
timestamp 1018054153
transform 1 0 5536 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8106
timestamp 1018054153
transform 1 0 5552 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8108
timestamp 1018054153
transform 1 0 5568 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8110
timestamp 1018054153
transform 1 0 5584 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8112
timestamp 1018054153
transform 1 0 5600 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8114
timestamp 1018054153
transform 1 0 5616 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8116
timestamp 1018054153
transform 1 0 5632 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8118
timestamp 1018054153
transform 1 0 5648 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8120
timestamp 1018054153
transform 1 0 5664 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8122
timestamp 1018054153
transform 1 0 5680 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8124
timestamp 1018054153
transform 1 0 5696 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8126
timestamp 1018054153
transform 1 0 5712 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8128
timestamp 1018054153
transform 1 0 5728 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8130
timestamp 1018054153
transform 1 0 5744 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8132
timestamp 1018054153
transform 1 0 5760 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8134
timestamp 1018054153
transform 1 0 5776 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8136
timestamp 1018054153
transform 1 0 5792 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8138
timestamp 1018054153
transform 1 0 5808 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8140
timestamp 1018054153
transform 1 0 5824 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8142
timestamp 1018054153
transform 1 0 5840 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8144
timestamp 1018054153
transform 1 0 5856 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8146
timestamp 1018054153
transform 1 0 5872 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8148
timestamp 1018054153
transform 1 0 5888 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8150
timestamp 1018054153
transform 1 0 5904 0 -1 2480
box -16 -6 32 210
use M2_M1  M2_M1_290
timestamp 1542725905
transform 1 0 5944 0 1 2310
box -4 -4 4 4
use FILL  FILL_8152
timestamp 1018054153
transform 1 0 5920 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8154
timestamp 1018054153
transform 1 0 5936 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8156
timestamp 1018054153
transform 1 0 5952 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8158
timestamp 1018054153
transform 1 0 5968 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8160
timestamp 1018054153
transform 1 0 5984 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8162
timestamp 1018054153
transform 1 0 6000 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8164
timestamp 1018054153
transform 1 0 6016 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8166
timestamp 1018054153
transform 1 0 6032 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8168
timestamp 1018054153
transform 1 0 6048 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8170
timestamp 1018054153
transform 1 0 6064 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8172
timestamp 1018054153
transform 1 0 6080 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8174
timestamp 1018054153
transform 1 0 6096 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8176
timestamp 1018054153
transform 1 0 6112 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8178
timestamp 1018054153
transform 1 0 6128 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8180
timestamp 1018054153
transform 1 0 6144 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8182
timestamp 1018054153
transform 1 0 6160 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8184
timestamp 1018054153
transform 1 0 6176 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8186
timestamp 1018054153
transform 1 0 6192 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8188
timestamp 1018054153
transform 1 0 6208 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8190
timestamp 1018054153
transform 1 0 6224 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8192
timestamp 1018054153
transform 1 0 6240 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8194
timestamp 1018054153
transform 1 0 6256 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8196
timestamp 1018054153
transform 1 0 6272 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8198
timestamp 1018054153
transform 1 0 6288 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8200
timestamp 1018054153
transform 1 0 6304 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8202
timestamp 1018054153
transform 1 0 6320 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8204
timestamp 1018054153
transform 1 0 6336 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8206
timestamp 1018054153
transform 1 0 6352 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8208
timestamp 1018054153
transform 1 0 6368 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8210
timestamp 1018054153
transform 1 0 6384 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8212
timestamp 1018054153
transform 1 0 6400 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8214
timestamp 1018054153
transform 1 0 6416 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8216
timestamp 1018054153
transform 1 0 6432 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8218
timestamp 1018054153
transform 1 0 6448 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8220
timestamp 1018054153
transform 1 0 6464 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8222
timestamp 1018054153
transform 1 0 6480 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8224
timestamp 1018054153
transform 1 0 6496 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8226
timestamp 1018054153
transform 1 0 6512 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8228
timestamp 1018054153
transform 1 0 6528 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8230
timestamp 1018054153
transform 1 0 6544 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8232
timestamp 1018054153
transform 1 0 6560 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8234
timestamp 1018054153
transform 1 0 6576 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8236
timestamp 1018054153
transform 1 0 6592 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8238
timestamp 1018054153
transform 1 0 6608 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8240
timestamp 1018054153
transform 1 0 6624 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8242
timestamp 1018054153
transform 1 0 6640 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8244
timestamp 1018054153
transform 1 0 6656 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8246
timestamp 1018054153
transform 1 0 6672 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8248
timestamp 1018054153
transform 1 0 6688 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8250
timestamp 1018054153
transform 1 0 6704 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8252
timestamp 1018054153
transform 1 0 6720 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8254
timestamp 1018054153
transform 1 0 6736 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8256
timestamp 1018054153
transform 1 0 6752 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8258
timestamp 1018054153
transform 1 0 6768 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8260
timestamp 1018054153
transform 1 0 6784 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8262
timestamp 1018054153
transform 1 0 6800 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8264
timestamp 1018054153
transform 1 0 6816 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8266
timestamp 1018054153
transform 1 0 6832 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8268
timestamp 1018054153
transform 1 0 6848 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8270
timestamp 1018054153
transform 1 0 6864 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8272
timestamp 1018054153
transform 1 0 6880 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8274
timestamp 1018054153
transform 1 0 6896 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8276
timestamp 1018054153
transform 1 0 6912 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8278
timestamp 1018054153
transform 1 0 6928 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8280
timestamp 1018054153
transform 1 0 6944 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8282
timestamp 1018054153
transform 1 0 6960 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8284
timestamp 1018054153
transform 1 0 6976 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8286
timestamp 1018054153
transform 1 0 6992 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8288
timestamp 1018054153
transform 1 0 7008 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8290
timestamp 1018054153
transform 1 0 7024 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8292
timestamp 1018054153
transform 1 0 7040 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8294
timestamp 1018054153
transform 1 0 7056 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8296
timestamp 1018054153
transform 1 0 7072 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8298
timestamp 1018054153
transform 1 0 7088 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8300
timestamp 1018054153
transform 1 0 7104 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8302
timestamp 1018054153
transform 1 0 7120 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8304
timestamp 1018054153
transform 1 0 7136 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8306
timestamp 1018054153
transform 1 0 7152 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8308
timestamp 1018054153
transform 1 0 7168 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8310
timestamp 1018054153
transform 1 0 7184 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8312
timestamp 1018054153
transform 1 0 7200 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8314
timestamp 1018054153
transform 1 0 7216 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8316
timestamp 1018054153
transform 1 0 7232 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8318
timestamp 1018054153
transform 1 0 7248 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8320
timestamp 1018054153
transform 1 0 7264 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8322
timestamp 1018054153
transform 1 0 7280 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8324
timestamp 1018054153
transform 1 0 7296 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8326
timestamp 1018054153
transform 1 0 7312 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8328
timestamp 1018054153
transform 1 0 7328 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8330
timestamp 1018054153
transform 1 0 7344 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8332
timestamp 1018054153
transform 1 0 7360 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8334
timestamp 1018054153
transform 1 0 7376 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8336
timestamp 1018054153
transform 1 0 7392 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8338
timestamp 1018054153
transform 1 0 7408 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8340
timestamp 1018054153
transform 1 0 7424 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8342
timestamp 1018054153
transform 1 0 7440 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8344
timestamp 1018054153
transform 1 0 7456 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8346
timestamp 1018054153
transform 1 0 7472 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8348
timestamp 1018054153
transform 1 0 7488 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8350
timestamp 1018054153
transform 1 0 7504 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8352
timestamp 1018054153
transform 1 0 7520 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8354
timestamp 1018054153
transform 1 0 7536 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8356
timestamp 1018054153
transform 1 0 7552 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8358
timestamp 1018054153
transform 1 0 7568 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8360
timestamp 1018054153
transform 1 0 7584 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8362
timestamp 1018054153
transform 1 0 7600 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8364
timestamp 1018054153
transform 1 0 7616 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8366
timestamp 1018054153
transform 1 0 7632 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8368
timestamp 1018054153
transform 1 0 7648 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8370
timestamp 1018054153
transform 1 0 7664 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8372
timestamp 1018054153
transform 1 0 7680 0 -1 2480
box -16 -6 32 210
use FILL  FILL_8374
timestamp 1018054153
transform 1 0 7696 0 -1 2480
box -16 -6 32 210
use M2_M1  M2_M1_291
timestamp 1542725905
transform 1 0 7848 0 1 2310
box -4 -4 4 4
use mult_pad_VIA1  mult_pad_VIA1_51
timestamp 1542725905
transform 1 0 7788 0 1 2280
box -48 -6 48 6
use FILL  FILL_8376
timestamp 1018054153
transform 1 0 7712 0 -1 2480
box -16 -6 32 210
use mult_pad_VIA0  mult_pad_VIA0_4
timestamp 1542725905
transform 1 0 2212 0 1 2220
box -48 -48 48 48
use mult_pad_VIA0  mult_pad_VIA0_5
timestamp 1542725905
transform 1 0 7788 0 1 2220
box -48 -48 48 48
use mult_pad_VIA0  mult_pad_VIA0_6
timestamp 1542725905
transform 1 0 2092 0 1 2100
box -48 -48 48 48
use M3_M2  M3_M2_128
timestamp 1542725905
transform 1 0 6520 0 1 2150
box -6 -6 6 6
use M3_M2  M3_M2_129
timestamp 1542725905
transform 1 0 6680 0 1 2150
box -6 -6 6 6
use mult_pad_VIA0  mult_pad_VIA0_7
timestamp 1542725905
transform 1 0 7908 0 1 2100
box -48 -48 48 48
use M2_M1  M2_M1_292
timestamp 1542725905
transform 1 0 7688 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_293
timestamp 1542725905
transform 1 0 7880 0 1 2030
box -4 -4 4 4
use PADNC  PADNC_9
timestamp 1084294400
transform 0 -1 2000 1 0 2000
box -6 -6 606 2000
use PADFC  PADFC_3
timestamp 949001400
transform 0 -1 2000 1 0 0
box 654 -6 2006 1346
use PADNC  PADNC_10
timestamp 1084294400
transform -1 0 2600 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_11
timestamp 1084294400
transform -1 0 3200 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_12
timestamp 1084294400
transform -1 0 3800 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_13
timestamp 1084294400
transform -1 0 4400 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_14
timestamp 1084294400
transform -1 0 5000 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_15
timestamp 1084294400
transform -1 0 5600 0 -1 2000
box -6 -6 606 2000
use PADNC  PADNC_16
timestamp 1084294400
transform -1 0 6200 0 -1 2000
box -6 -6 606 2000
use PADOUT  PADOUT_6
timestamp 1084294529
transform -1 0 6800 0 -1 2000
box -12 -6 606 2000
use PADOUT  PADOUT_7
timestamp 1084294529
transform -1 0 7400 0 -1 2000
box -12 -6 606 2000
use PADOUT  PADOUT_5
timestamp 1084294529
transform 0 1 8000 -1 0 2600
box -12 -6 606 2000
use PADFC  PADFC_2
timestamp 949001400
transform -1 0 10000 0 -1 2000
box 654 -6 2006 1346
use PADOUT  PADOUT_8
timestamp 1084294529
transform -1 0 8000 0 -1 2000
box -12 -6 606 2000
<< labels >>
rlabel metal3 7116 264 7116 264 4 result[7]
rlabel metal3 7716 264 7716 264 4 result[6]
rlabel metal3 9736 2316 9736 2316 4 result[5]
rlabel metal3 9736 2916 9736 2916 4 result[4]
rlabel metal3 9736 3516 9736 3516 4 result[3]
rlabel metal3 9736 4116 9736 4116 4 result[2]
rlabel metal3 9736 4716 9736 4716 4 result[1]
rlabel metal3 9736 5316 9736 5316 4 result[0]
rlabel metal3 6516 264 6516 264 4 cout
rlabel metal3 4692 9762 4692 9762 4 a[3]
rlabel metal3 5292 9762 5292 9762 4 a[2]
rlabel metal3 5892 9762 5892 9762 4 a[1]
rlabel metal3 6492 9762 6492 9762 4 a[0]
rlabel metal3 238 3492 238 3492 4 b[3]
rlabel metal3 238 4092 238 4092 4 b[2]
rlabel metal3 238 4692 238 4692 4 b[1]
rlabel metal3 238 5292 238 5292 4 b[0]
rlabel metal3 238 5892 238 5892 4 reset
rlabel metal3 238 6492 238 6492 4 clk
rlabel metal2 2044 2052 2044 2052 4 gnd
rlabel metal2 2164 2172 2164 2172 4 vdd
rlabel metal3 9672 7662 9678 7670 0 gnd
rlabel metal3 9684 7016 9684 7018 0 vdd
rlabel metal3 202 7192 204 7192 0 vdd
rlabel metal3 220 7748 226 7748 0 gnd
<< end >>
