* SPICE3 file created from bs2.ext - technology: scmos

.option scale=0.3u

M1000 dffpos_0/a_35_65# dffpos_0/clk_b gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=540 ps=298
M1001 dffpos_0/clk dffpos_0/clk_b dffpos_0/a_35_65# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1002 dffpos_0/a_56_65# dffpos_0/D gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1003 dffpos_0/a_61_9# dffpos_0/clk_b dffpos_0/a_56_65# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1004 dffpos_0/a_69_65# dffpos_0/clk dffpos_0/a_61_9# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1005 gnd dffpos_0/a_72_7# dffpos_0/a_69_65# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 dffpos_0/a_72_7# dffpos_0/a_61_9# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1007 dffpos_0/a_99_65# dffpos_0/a_72_7# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1008 dffpos_0/a_104_9# dffpos_0/clk dffpos_0/a_99_65# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1009 dffpos_0/a_112_65# dffpos_0/clk_b dffpos_0/a_104_9# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1010 gnd Out dffpos_0/a_112_65# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 dffpos_0/a_126_65# dffpos_0/a_104_9# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1012 Out dffpos_0/a_104_9# dffpos_0/a_126_65# Gnd nfet w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1013 dffpos_0/a_35_9# dffpos_0/clk_b vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=980 ps=458
M1014 dffpos_0/clk dffpos_0/clk_b dffpos_0/a_35_9# Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 dffpos_0/a_56_9# dffpos_0/D vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1016 dffpos_0/a_61_9# dffpos_0/clk dffpos_0/a_56_9# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1017 dffpos_0/a_69_9# dffpos_0/clk_b dffpos_0/a_61_9# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1018 vdd dffpos_0/a_72_7# dffpos_0/a_69_9# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 dffpos_0/a_72_7# dffpos_0/a_61_9# vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1020 dffpos_0/a_99_9# dffpos_0/a_72_7# vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1021 dffpos_0/a_104_9# dffpos_0/clk_b dffpos_0/a_99_9# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1022 dffpos_0/a_112_9# dffpos_0/clk dffpos_0/a_104_9# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1023 vdd Out dffpos_0/a_112_9# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 dffpos_0/a_126_9# dffpos_0/a_104_9# vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1025 Out dffpos_0/a_104_9# dffpos_0/a_126_9# Vdd pfet w=20 l=2
+  ad=150 pd=80 as=0 ps=0
M1026 dffpos_0/clk_b en vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1027 vdd clk dffpos_0/clk_b Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 nand_0/a_9_6# en gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1029 dffpos_0/clk_b clk nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1030 bc1a_0/inverter_1/Y Init vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1031 bc1a_0/inverter_1/Y Init gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1032 muxB_in Init Out Vdd pfet w=10 l=2
+  ad=110 pd=62 as=0 ps=0
M1033 mplier bc1a_0/inverter_1/Y muxB_in Vdd pfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 muxB_in bc1a_0/inverter_1/Y Out Gnd nfet w=10 l=2
+  ad=110 pd=62 as=0 ps=0
M1035 mplier Init muxB_in Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1036 dffpos_0/D bc1a_0/inverter_1/Y muxA_in Gnd nfet w=10 l=2
+  ad=60 pd=32 as=50 ps=30
M1037 muxB_in Init dffpos_0/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 dffpos_0/D Init muxA_in Vdd pfet w=10 l=2
+  ad=60 pd=32 as=50 ps=30
M1039 muxB_in bc1a_0/inverter_1/Y dffpos_0/D Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 a_52_99# q0 vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1041 muxA_out q0 gnd Vdd pfet w=10 l=2
+  ad=60 pd=32 as=466 ps=446
M1042 mcand a_52_99# muxA_out Vdd pfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1043 muxA_out a_52_99# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1044 mcand q0 muxA_out Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1045 a_52_99# q0 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 muxA_out gnd 2.296470fF
C1 dffpos_0/clk dffpos_0/D 2.254440fF
C2 mcand gnd! 8.794080fF
C3 muxA_out gnd! 4.703610fF
C4 a_52_99# gnd! 7.399800fF
C5 q0 gnd! 12.861000fF
C6 clk gnd! 10.136520fF
C7 vdd gnd! 53.604695fF
C8 muxA_in gnd! 9.437399fF
C9 mplier gnd! 2.239920fF
C10 muxB_in gnd! 12.985920fF
C11 Init gnd! 13.238681fF
C12 bc1a_0/inverter_1/Y gnd! 11.778479fF
C13 en gnd! 10.362309fF
C14 dffpos_0/a_104_9# gnd! 4.015080fF
C15 Out gnd! 12.704761fF
C16 dffpos_0/a_61_9# gnd! 3.452040fF
C17 dffpos_0/a_72_7# gnd! 4.794840fF
C18 dffpos_0/clk gnd! 7.541550fF
C19 dffpos_0/D gnd! 6.984990fF
C20 dffpos_0/clk_b gnd! 9.353609fF
C21 gnd gnd! 43.963902fF
