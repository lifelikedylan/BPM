magic
tech scmos
timestamp 1542725905
<< metal1 >>
rect -2 2 2 3
rect -2 -3 2 -2
<< m2contact >>
rect -2 -2 2 2
<< metal2 >>
rect -2 2 2 3
rect -2 -3 2 -2
<< end >>
