magic
tech scmos
timestamp 1543282957
use ../../bs1/magic/bs1  bs1_0 ../../bs1/magic
array 0 0 220 0 7 180
timestamp 1543282590
transform 1 0 1 0 1 3
box -2 -3 218 177
<< end >>
