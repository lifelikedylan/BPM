magic
tech scmos
timestamp 1543281763
<< ntransistor >>
rect -18 -18 -16 -8
rect -10 -18 -8 -8
<< ptransistor >>
rect -18 24 -16 34
rect -10 24 -8 34
<< ndiffusion >>
rect -19 -18 -18 -8
rect -16 -18 -15 -8
rect -11 -18 -10 -8
rect -8 -18 -7 -8
<< pdiffusion >>
rect -19 24 -18 34
rect -16 24 -15 34
rect -11 24 -10 34
rect -8 24 -7 34
<< ndcontact >>
rect -23 -18 -19 -8
rect -15 -18 -11 -8
rect -7 -18 -3 -8
<< pdcontact >>
rect -23 24 -19 34
rect -15 24 -11 34
rect -7 24 -3 34
<< psubstratepcontact >>
rect -23 -36 -19 -32
rect -7 -36 -3 -32
<< nsubstratencontact >>
rect -25 42 -21 46
rect -6 42 -2 46
<< polysilicon >>
rect -26 35 -16 37
rect -18 34 -16 35
rect -10 34 -8 36
rect -18 -1 -16 24
rect -10 23 -8 24
rect -10 21 0 23
rect -18 -3 -8 -1
rect -18 -8 -16 -6
rect -10 -8 -8 -3
rect -18 -23 -16 -18
rect -10 -20 -8 -18
rect -18 -25 0 -23
<< polycontact >>
rect -30 34 -26 38
rect 0 20 4 24
rect 0 -26 4 -22
<< metal1 >>
rect -30 46 4 47
rect -30 42 -25 46
rect -21 42 -6 46
rect -2 42 4 46
rect -30 41 4 42
rect -30 11 -26 34
rect -23 -8 -19 24
rect -15 -8 -11 24
rect -7 -8 -3 24
rect -23 -24 -19 -18
rect -30 -28 -19 -24
rect 0 -22 4 20
rect -30 -32 4 -31
rect -30 -36 -23 -32
rect -19 -36 -7 -32
rect -3 -36 4 -32
rect -30 -37 4 -36
<< labels >>
rlabel polycontact 2 22 2 22 0 Sel_bar
rlabel polycontact -28 36 -28 36 0 Sel
rlabel nsubstratencontact -3 43 -3 43 3 Vdd
rlabel metal1 -28 -26 -28 -26 3 In_0
rlabel metal1 -5 10 -5 11 1 in_1
rlabel metal1 -13 15 -13 15 3 Out
<< end >>
