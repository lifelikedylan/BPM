VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rca8
  CLASS RING ;
  ORIGIN 4.8 4.8 ;
  FOREIGN rca8 -4.8 -4.8 ;
  SIZE 278.4 BY 48.3 ;
  SYMMETRY X Y R90 ;
  PIN a_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12 36.6 13.2 38.7 ;
    END
  END a_0
  PIN a_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 54 36.6 55.2 38.7 ;
    END
  END a_1
  PIN a_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 79.2 36.6 80.4 38.7 ;
    END
  END a_2
  PIN a_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 121.2 36.6 122.4 38.7 ;
    END
  END a_3
  PIN a_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 146.4 36.6 147.6 38.7 ;
    END
  END a_4
  PIN a_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 188.4 36.6 189.6 38.7 ;
    END
  END a_5
  PIN a_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 213.6 36.6 214.8 38.7 ;
    END
  END a_6
  PIN a_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 255.6 36.6 256.8 38.7 ;
    END
  END a_7
  PIN b_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15 34.2 16.2 38.7 ;
    END
  END b_0
  PIN b_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51 34.2 52.2 38.7 ;
    END
  END b_1
  PIN b_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 82.2 34.2 83.4 38.7 ;
    END
  END b_2
  PIN b_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 118.2 34.2 119.4 38.7 ;
    END
  END b_3
  PIN b_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 149.4 34.2 150.6 38.7 ;
    END
  END b_4
  PIN b_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 185.4 34.2 186.6 38.7 ;
    END
  END b_5
  PIN b_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 216.6 34.2 217.8 38.7 ;
    END
  END b_6
  PIN b_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 252.6 34.2 253.8 38.7 ;
    END
  END b_7
  PIN c_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18 31.8 19.2 38.7 ;
    END
  END c_0
  PIN cout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 255.6 0 256.8 1.8 ;
    END
  END cout
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER metal1 ;
        RECT 265.8 0.6 268.8 38.7 ;
        RECT 198.6 37.8 204.6 38.7 ;
        RECT 131.4 37.8 137.4 38.7 ;
        RECT 64.2 37.8 70.2 38.7 ;
        RECT 0 0.6 3 38.7 ;
    END
  END gnd
  PIN sum_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15 0 16.2 0.6 ;
    END
  END sum_0
  PIN sum_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51 0 52.2 0.6 ;
    END
  END sum_1
  PIN sum_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 82.2 0 83.4 0.6 ;
    END
  END sum_2
  PIN sum_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 118.2 0 119.4 0.6 ;
    END
  END sum_3
  PIN sum_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 149.4 0 150.6 0.6 ;
    END
  END sum_4
  PIN sum_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 185.4 0 186.6 0.6 ;
    END
  END sum_5
  PIN sum_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 216.6 0 217.8 0.6 ;
    END
  END sum_6
  PIN sum_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 252.6 0 253.8 0.6 ;
    END
  END sum_7
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER metal1 ;
        RECT 232.8 37.8 237.6 38.7 ;
        RECT 234.6 0.6 235.8 38.7 ;
        RECT 165.6 37.8 170.4 38.7 ;
        RECT 98.4 37.8 103.2 38.7 ;
        RECT 31.2 38.1 36 38.7 ;
        RECT 33 0.6 34.2 38.7 ;
    END
  END vdd
  OBS
    LAYER metal2 ;
      RECT 260.7 1.8 261.9 3 ;
      RECT 255.6 1.8 256.8 3 ;
      RECT 244.5 1.8 245.7 3 ;
      RECT 244.5 1.8 261.9 2.7 ;
      RECT 258 28.2 261.9 29.4 ;
      RECT 244.5 28.2 248.1 29.4 ;
      RECT 244.5 28.2 261.9 29.1 ;
      RECT 252.6 6.6 253.8 7.8 ;
      RECT 244.5 6.6 245.7 7.8 ;
      RECT 244.5 6.6 261 7.5 ;
      RECT 259.8 6 261 7.5 ;
      RECT 231 30.9 250.8 31.8 ;
      RECT 249.6 30.6 250.8 31.8 ;
      RECT 231 1.8 231.9 31.8 ;
      RECT 224.7 1.8 225.9 3 ;
      RECT 213.6 1.8 214.8 3 ;
      RECT 208.5 1.8 209.7 3 ;
      RECT 208.5 1.8 231.9 2.7 ;
      RECT 224.7 6.6 225.9 7.8 ;
      RECT 216.6 6.6 217.8 7.8 ;
      RECT 209.4 6.6 225.9 7.5 ;
      RECT 209.4 6 210.6 7.5 ;
      RECT 222.3 28.2 225.9 29.4 ;
      RECT 208.5 28.2 212.4 29.4 ;
      RECT 208.5 28.2 225.9 29.1 ;
      RECT 196.5 30.9 220.8 31.8 ;
      RECT 219.6 30.6 220.8 31.8 ;
      RECT 196.5 1.8 197.7 31.8 ;
      RECT 193.5 1.8 194.7 3 ;
      RECT 188.4 1.8 189.6 3 ;
      RECT 177.3 1.8 178.5 3 ;
      RECT 177.3 1.8 197.7 2.7 ;
      RECT 190.8 28.2 194.7 29.4 ;
      RECT 177.3 28.2 180.9 29.4 ;
      RECT 177.3 28.2 194.7 29.1 ;
      RECT 185.4 6.6 186.6 7.8 ;
      RECT 177.3 6.6 178.5 7.8 ;
      RECT 177.3 6.6 193.8 7.5 ;
      RECT 192.6 6 193.8 7.5 ;
      RECT 163.8 30.9 183.6 31.8 ;
      RECT 182.4 30.6 183.6 31.8 ;
      RECT 163.8 1.8 164.7 31.8 ;
      RECT 157.5 1.8 158.7 3 ;
      RECT 146.4 1.8 147.6 3 ;
      RECT 141.3 1.8 142.5 3 ;
      RECT 141.3 1.8 164.7 2.7 ;
      RECT 157.5 6.6 158.7 7.8 ;
      RECT 149.4 6.6 150.6 7.8 ;
      RECT 142.2 6.6 158.7 7.5 ;
      RECT 142.2 6 143.4 7.5 ;
      RECT 155.1 28.2 158.7 29.4 ;
      RECT 141.3 28.2 145.2 29.4 ;
      RECT 141.3 28.2 158.7 29.1 ;
      RECT 152.4 30.6 153.6 31.8 ;
      RECT 129.6 30.6 153.6 31.5 ;
      RECT 129.6 1.8 130.5 31.5 ;
      RECT 126.3 1.8 127.5 3 ;
      RECT 121.2 1.8 122.4 3 ;
      RECT 110.1 1.8 111.3 3 ;
      RECT 110.1 1.8 130.5 2.7 ;
      RECT 123.6 28.2 127.5 29.4 ;
      RECT 110.1 28.2 113.7 29.4 ;
      RECT 110.1 28.2 127.5 29.1 ;
      RECT 118.2 6.6 119.4 7.8 ;
      RECT 110.1 6.6 111.3 7.8 ;
      RECT 110.1 6.6 126.6 7.5 ;
      RECT 125.4 6 126.6 7.5 ;
      RECT 96.6 30.9 116.4 31.8 ;
      RECT 115.2 30.6 116.4 31.8 ;
      RECT 96.6 1.8 97.5 31.8 ;
      RECT 90.3 1.8 91.5 3 ;
      RECT 79.2 1.8 80.4 3 ;
      RECT 74.1 1.8 75.3 3 ;
      RECT 74.1 1.8 97.5 2.7 ;
      RECT 90.3 6.6 91.5 7.8 ;
      RECT 82.2 6.6 83.4 7.8 ;
      RECT 75 6.6 91.5 7.5 ;
      RECT 75 6 76.2 7.5 ;
      RECT 87.9 28.2 91.5 29.4 ;
      RECT 74.1 28.2 78 29.4 ;
      RECT 74.1 28.2 91.5 29.1 ;
      RECT 62.4 30.9 86.4 31.8 ;
      RECT 85.2 30.6 86.4 31.8 ;
      RECT 62.4 1.8 63.3 31.8 ;
      RECT 59.1 1.8 60.3 3 ;
      RECT 54 1.8 55.2 3 ;
      RECT 42.9 1.8 44.1 3 ;
      RECT 42.9 1.8 63.3 2.7 ;
      RECT 56.4 28.2 60.3 29.4 ;
      RECT 42.9 28.2 46.5 29.4 ;
      RECT 42.9 28.2 60.3 29.1 ;
      RECT 51 6.6 52.2 7.8 ;
      RECT 42.9 6.6 44.1 7.8 ;
      RECT 42.9 6.6 59.4 7.5 ;
      RECT 58.2 6 59.4 7.5 ;
      RECT 29.4 30.9 49.2 31.8 ;
      RECT 48 30.6 49.2 31.8 ;
      RECT 29.4 1.8 30.3 31.8 ;
      RECT 23.1 1.8 24.3 3 ;
      RECT 12 1.8 13.2 3 ;
      RECT 6.9 1.8 8.1 3 ;
      RECT 6.9 1.8 30.3 2.7 ;
      RECT 23.1 6.6 24.3 7.8 ;
      RECT 15 6.6 16.2 7.8 ;
      RECT 7.8 6.6 24.3 7.5 ;
      RECT 7.8 6 9 7.5 ;
      RECT 20.7 28.2 24.3 29.4 ;
      RECT 6.9 28.2 10.8 29.4 ;
      RECT 6.9 28.2 24.3 29.1 ;
      RECT 243.6 13.8 261.9 15 ;
      RECT 208.5 13.8 226.8 15 ;
      RECT 176.4 13.8 194.7 15 ;
      RECT 141.3 13.8 159.6 15 ;
      RECT 109.2 13.8 127.5 15 ;
      RECT 74.1 13.8 92.4 15 ;
      RECT 42 13.8 60.3 15 ;
      RECT 6.9 13.8 25.2 15 ;
      RECT 18 30.6 19.2 31.8 ;
    LAYER metal1 ;
      RECT 261.9 6.6 264.9 7.8 ;
      RECT 259.8 6.3 262.8 7.2 ;
      RECT 259.8 6 261 7.2 ;
      RECT 261.9 14.4 264.9 15.9 ;
      RECT 260.7 13.8 261.9 15.3 ;
      RECT 259.8 8.1 260.7 14.7 ;
      RECT 259.8 8.1 261 9.3 ;
      RECT 261.9 21.9 264.9 23.1 ;
      RECT 260.1 21.9 264.9 22.8 ;
      RECT 260.1 17.4 261 22.8 ;
      RECT 260.1 17.4 264.9 18.3 ;
      RECT 261.9 17.1 264.9 18.3 ;
      RECT 261.9 35.4 264.9 36.6 ;
      RECT 260.1 35.4 264.9 36.3 ;
      RECT 260.1 30.9 261 36.3 ;
      RECT 260.1 30.9 264.9 31.8 ;
      RECT 261.9 30.6 264.9 31.8 ;
      RECT 258 28.2 259.2 29.4 ;
      RECT 258 5.1 258.9 29.4 ;
      RECT 258 15.9 259.2 17.1 ;
      RECT 257.7 5.1 258.9 6.3 ;
      RECT 255.6 33.9 256.8 35.7 ;
      RECT 255.9 9.6 256.8 35.7 ;
      RECT 255.6 23.1 256.8 24.3 ;
      RECT 255.6 9.6 256.8 10.8 ;
      RECT 252.6 31.5 253.8 33.3 ;
      RECT 252.6 11.7 253.5 33.3 ;
      RECT 252.3 26.7 253.5 27.9 ;
      RECT 252.6 20.7 253.8 21.9 ;
      RECT 252.3 11.7 253.5 12.9 ;
      RECT 249.6 29.1 250.8 31.8 ;
      RECT 249.6 13.8 250.5 31.8 ;
      RECT 249.6 18.3 250.8 19.5 ;
      RECT 249.6 13.8 250.8 15 ;
      RECT 246.9 28.2 248.1 29.4 ;
      RECT 247.2 5.1 248.1 29.4 ;
      RECT 247.2 15.9 248.4 17.1 ;
      RECT 246.9 5.1 248.1 6.3 ;
      RECT 238.5 21.9 244.5 23.1 ;
      RECT 238.5 21.9 246.3 22.8 ;
      RECT 245.4 17.4 246.3 22.8 ;
      RECT 238.5 17.4 246.3 18.3 ;
      RECT 238.5 17.1 244.5 18.3 ;
      RECT 238.5 35.4 244.5 36.6 ;
      RECT 238.5 35.4 246.3 36.3 ;
      RECT 245.4 30.9 246.3 36.3 ;
      RECT 238.5 30.9 246.3 31.8 ;
      RECT 238.5 30.6 244.5 31.8 ;
      RECT 238.5 14.4 244.5 15.9 ;
      RECT 243.6 13.8 245.7 15 ;
      RECT 236.7 0.6 237.6 36.9 ;
      RECT 236.7 33 244.5 34.2 ;
      RECT 236.7 24.3 244.5 25.5 ;
      RECT 236.7 19.5 244.5 20.7 ;
      RECT 236.7 9 244.5 10.2 ;
      RECT 236.7 4.2 244.5 5.4 ;
      RECT 232.8 0.6 233.7 36.9 ;
      RECT 225.9 33 233.7 34.2 ;
      RECT 225.9 24.3 233.7 25.5 ;
      RECT 225.9 19.5 233.7 20.7 ;
      RECT 225.9 9 233.7 10.2 ;
      RECT 225.9 4.2 233.7 5.4 ;
      RECT 225.9 14.4 231.9 15.9 ;
      RECT 224.7 13.8 226.8 15 ;
      RECT 225.9 21.9 231.9 23.1 ;
      RECT 224.1 21.9 231.9 22.8 ;
      RECT 224.1 17.4 225 22.8 ;
      RECT 224.1 17.4 231.9 18.3 ;
      RECT 225.9 17.1 231.9 18.3 ;
      RECT 225.9 35.4 231.9 36.6 ;
      RECT 224.1 35.4 231.9 36.3 ;
      RECT 224.1 30.9 225 36.3 ;
      RECT 224.1 30.9 231.9 31.8 ;
      RECT 225.9 30.6 231.9 31.8 ;
      RECT 222.3 28.2 223.5 29.4 ;
      RECT 222.3 5.1 223.2 29.4 ;
      RECT 222 15.9 223.2 17.1 ;
      RECT 222.3 5.1 223.5 6.3 ;
      RECT 219.6 29.1 220.8 31.8 ;
      RECT 219.9 13.8 220.8 31.8 ;
      RECT 219.6 18.3 220.8 19.5 ;
      RECT 219.6 13.8 220.8 15 ;
      RECT 216.6 31.5 217.8 33.3 ;
      RECT 216.9 11.7 217.8 33.3 ;
      RECT 216.9 26.7 218.1 27.9 ;
      RECT 216.6 20.7 217.8 21.9 ;
      RECT 216.9 11.7 218.1 12.9 ;
      RECT 213.6 33.9 214.8 35.7 ;
      RECT 213.6 9.6 214.5 35.7 ;
      RECT 213.6 23.1 214.8 24.3 ;
      RECT 213.6 9.6 214.8 10.8 ;
      RECT 211.2 28.2 212.4 29.4 ;
      RECT 211.5 5.1 212.4 29.4 ;
      RECT 211.2 15.9 212.4 17.1 ;
      RECT 211.5 5.1 212.7 6.3 ;
      RECT 205.5 6.6 208.5 7.8 ;
      RECT 209.4 6 210.6 7.2 ;
      RECT 207.6 6.3 210.6 7.2 ;
      RECT 205.5 14.4 208.5 15.9 ;
      RECT 205.5 14.4 209.7 15.3 ;
      RECT 209.7 8.1 210.6 14.7 ;
      RECT 208.5 13.8 210.6 14.7 ;
      RECT 209.4 8.1 210.6 9.3 ;
      RECT 205.5 21.9 208.5 23.1 ;
      RECT 205.5 21.9 210.3 22.8 ;
      RECT 209.4 17.4 210.3 22.8 ;
      RECT 205.5 17.4 210.3 18.3 ;
      RECT 205.5 17.1 208.5 18.3 ;
      RECT 205.5 35.4 208.5 36.6 ;
      RECT 205.5 35.4 210.3 36.3 ;
      RECT 209.4 30.9 210.3 36.3 ;
      RECT 205.5 30.9 210.3 31.8 ;
      RECT 205.5 30.6 208.5 31.8 ;
      RECT 198.6 0.6 204.6 36.9 ;
      RECT 194.7 33 208.5 34.2 ;
      RECT 194.7 24.3 208.5 25.5 ;
      RECT 194.7 19.5 208.5 20.7 ;
      RECT 194.7 9 208.5 10.2 ;
      RECT 194.7 4.2 208.5 5.4 ;
      RECT 194.7 6.6 197.7 7.8 ;
      RECT 192.6 6.3 195.6 7.2 ;
      RECT 192.6 6 193.8 7.2 ;
      RECT 194.7 14.4 197.7 15.9 ;
      RECT 193.5 13.8 194.7 15.3 ;
      RECT 192.6 8.1 193.5 14.7 ;
      RECT 192.6 8.1 193.8 9.3 ;
      RECT 194.7 21.9 197.7 23.1 ;
      RECT 192.9 21.9 197.7 22.8 ;
      RECT 192.9 17.4 193.8 22.8 ;
      RECT 192.9 17.4 197.7 18.3 ;
      RECT 194.7 17.1 197.7 18.3 ;
      RECT 194.7 35.4 197.7 36.6 ;
      RECT 192.9 35.4 197.7 36.3 ;
      RECT 192.9 30.9 193.8 36.3 ;
      RECT 192.9 30.9 197.7 31.8 ;
      RECT 194.7 30.6 197.7 31.8 ;
      RECT 190.8 28.2 192 29.4 ;
      RECT 190.8 5.1 191.7 29.4 ;
      RECT 190.8 15.9 192 17.1 ;
      RECT 190.5 5.1 191.7 6.3 ;
      RECT 188.4 33.9 189.6 35.7 ;
      RECT 188.7 9.6 189.6 35.7 ;
      RECT 188.4 23.1 189.6 24.3 ;
      RECT 188.4 9.6 189.6 10.8 ;
      RECT 185.4 31.5 186.6 33.3 ;
      RECT 185.4 11.7 186.3 33.3 ;
      RECT 185.1 26.7 186.3 27.9 ;
      RECT 185.4 20.7 186.6 21.9 ;
      RECT 185.1 11.7 186.3 12.9 ;
      RECT 182.4 29.1 183.6 31.8 ;
      RECT 182.4 13.8 183.3 31.8 ;
      RECT 182.4 18.3 183.6 19.5 ;
      RECT 182.4 13.8 183.6 15 ;
      RECT 179.7 28.2 180.9 29.4 ;
      RECT 180 5.1 180.9 29.4 ;
      RECT 180 15.9 181.2 17.1 ;
      RECT 179.7 5.1 180.9 6.3 ;
      RECT 171.3 21.9 177.3 23.1 ;
      RECT 171.3 21.9 179.1 22.8 ;
      RECT 178.2 17.4 179.1 22.8 ;
      RECT 171.3 17.4 179.1 18.3 ;
      RECT 171.3 17.1 177.3 18.3 ;
      RECT 171.3 35.4 177.3 36.6 ;
      RECT 171.3 35.4 179.1 36.3 ;
      RECT 178.2 30.9 179.1 36.3 ;
      RECT 171.3 30.9 179.1 31.8 ;
      RECT 171.3 30.6 177.3 31.8 ;
      RECT 171.3 14.4 177.3 15.9 ;
      RECT 176.4 13.8 178.5 15 ;
      RECT 165.6 0.6 170.4 36.9 ;
      RECT 158.7 33 177.3 34.2 ;
      RECT 158.7 24.3 177.3 25.5 ;
      RECT 158.7 19.5 177.3 20.7 ;
      RECT 158.7 9 177.3 10.2 ;
      RECT 158.7 4.2 177.3 5.4 ;
      RECT 158.7 14.4 164.7 15.9 ;
      RECT 157.5 13.8 159.6 15 ;
      RECT 158.7 21.9 164.7 23.1 ;
      RECT 156.9 21.9 164.7 22.8 ;
      RECT 156.9 17.4 157.8 22.8 ;
      RECT 156.9 17.4 164.7 18.3 ;
      RECT 158.7 17.1 164.7 18.3 ;
      RECT 158.7 35.4 164.7 36.6 ;
      RECT 156.9 35.4 164.7 36.3 ;
      RECT 156.9 30.9 157.8 36.3 ;
      RECT 156.9 30.9 164.7 31.8 ;
      RECT 158.7 30.6 164.7 31.8 ;
      RECT 155.1 28.2 156.3 29.4 ;
      RECT 155.1 5.1 156 29.4 ;
      RECT 154.8 15.9 156 17.1 ;
      RECT 155.1 5.1 156.3 6.3 ;
      RECT 152.4 29.1 153.6 31.8 ;
      RECT 152.7 13.8 153.6 31.8 ;
      RECT 152.4 18.3 153.6 19.5 ;
      RECT 152.4 13.8 153.6 15 ;
      RECT 149.4 31.5 150.6 33.3 ;
      RECT 149.7 11.7 150.6 33.3 ;
      RECT 149.7 26.7 150.9 27.9 ;
      RECT 149.4 20.7 150.6 21.9 ;
      RECT 149.7 11.7 150.9 12.9 ;
      RECT 146.4 33.9 147.6 35.7 ;
      RECT 146.4 9.6 147.3 35.7 ;
      RECT 146.4 23.1 147.6 24.3 ;
      RECT 146.4 9.6 147.6 10.8 ;
      RECT 144 28.2 145.2 29.4 ;
      RECT 144.3 5.1 145.2 29.4 ;
      RECT 144 15.9 145.2 17.1 ;
      RECT 144.3 5.1 145.5 6.3 ;
      RECT 138.3 6.6 141.3 7.8 ;
      RECT 142.2 6 143.4 7.2 ;
      RECT 140.4 6.3 143.4 7.2 ;
      RECT 138.3 14.4 141.3 15.9 ;
      RECT 138.3 14.4 142.5 15.3 ;
      RECT 142.5 8.1 143.4 14.7 ;
      RECT 141.3 13.8 143.4 14.7 ;
      RECT 142.2 8.1 143.4 9.3 ;
      RECT 138.3 21.9 141.3 23.1 ;
      RECT 138.3 21.9 143.1 22.8 ;
      RECT 142.2 17.4 143.1 22.8 ;
      RECT 138.3 17.4 143.1 18.3 ;
      RECT 138.3 17.1 141.3 18.3 ;
      RECT 138.3 35.4 141.3 36.6 ;
      RECT 138.3 35.4 143.1 36.3 ;
      RECT 142.2 30.9 143.1 36.3 ;
      RECT 138.3 30.9 143.1 31.8 ;
      RECT 138.3 30.6 141.3 31.8 ;
      RECT 131.4 0.6 137.4 36.9 ;
      RECT 127.5 33 141.3 34.2 ;
      RECT 127.5 24.3 141.3 25.5 ;
      RECT 127.5 19.5 141.3 20.7 ;
      RECT 127.5 9 141.3 10.2 ;
      RECT 127.5 4.2 141.3 5.4 ;
      RECT 127.5 6.6 130.5 7.8 ;
      RECT 125.4 6.3 128.4 7.2 ;
      RECT 125.4 6 126.6 7.2 ;
      RECT 127.5 14.4 130.5 15.9 ;
      RECT 126.3 13.8 127.5 15.3 ;
      RECT 125.4 8.1 126.3 14.7 ;
      RECT 125.4 8.1 126.6 9.3 ;
      RECT 127.5 21.9 130.5 23.1 ;
      RECT 125.7 21.9 130.5 22.8 ;
      RECT 125.7 17.4 126.6 22.8 ;
      RECT 125.7 17.4 130.5 18.3 ;
      RECT 127.5 17.1 130.5 18.3 ;
      RECT 127.5 35.4 130.5 36.6 ;
      RECT 125.7 35.4 130.5 36.3 ;
      RECT 125.7 30.9 126.6 36.3 ;
      RECT 125.7 30.9 130.5 31.8 ;
      RECT 127.5 30.6 130.5 31.8 ;
      RECT 123.6 28.2 124.8 29.4 ;
      RECT 123.6 5.1 124.5 29.4 ;
      RECT 123.6 15.9 124.8 17.1 ;
      RECT 123.3 5.1 124.5 6.3 ;
      RECT 121.2 33.9 122.4 35.7 ;
      RECT 121.5 9.6 122.4 35.7 ;
      RECT 121.2 23.1 122.4 24.3 ;
      RECT 121.2 9.6 122.4 10.8 ;
      RECT 118.2 31.5 119.4 33.3 ;
      RECT 118.2 11.7 119.1 33.3 ;
      RECT 117.9 26.7 119.1 27.9 ;
      RECT 118.2 20.7 119.4 21.9 ;
      RECT 117.9 11.7 119.1 12.9 ;
      RECT 115.2 29.1 116.4 31.8 ;
      RECT 115.2 13.8 116.1 31.8 ;
      RECT 115.2 18.3 116.4 19.5 ;
      RECT 115.2 13.8 116.4 15 ;
      RECT 112.5 28.2 113.7 29.4 ;
      RECT 112.8 5.1 113.7 29.4 ;
      RECT 112.8 15.9 114 17.1 ;
      RECT 112.5 5.1 113.7 6.3 ;
      RECT 104.1 21.9 110.1 23.1 ;
      RECT 104.1 21.9 111.9 22.8 ;
      RECT 111 17.4 111.9 22.8 ;
      RECT 104.1 17.4 111.9 18.3 ;
      RECT 104.1 17.1 110.1 18.3 ;
      RECT 104.1 35.4 110.1 36.6 ;
      RECT 104.1 35.4 111.9 36.3 ;
      RECT 111 30.9 111.9 36.3 ;
      RECT 104.1 30.9 111.9 31.8 ;
      RECT 104.1 30.6 110.1 31.8 ;
      RECT 104.1 14.4 110.1 15.9 ;
      RECT 109.2 13.8 111.3 15 ;
      RECT 98.4 0.6 103.2 36.9 ;
      RECT 91.5 33 110.1 34.2 ;
      RECT 91.5 24.3 110.1 25.5 ;
      RECT 91.5 19.5 110.1 20.7 ;
      RECT 91.5 9 110.1 10.2 ;
      RECT 91.5 4.2 110.1 5.4 ;
      RECT 91.5 14.4 97.5 15.9 ;
      RECT 90.3 13.8 92.4 15 ;
      RECT 91.5 21.9 97.5 23.1 ;
      RECT 89.7 21.9 97.5 22.8 ;
      RECT 89.7 17.4 90.6 22.8 ;
      RECT 89.7 17.4 97.5 18.3 ;
      RECT 91.5 17.1 97.5 18.3 ;
      RECT 91.5 35.4 97.5 36.6 ;
      RECT 89.7 35.4 97.5 36.3 ;
      RECT 89.7 30.9 90.6 36.3 ;
      RECT 89.7 30.9 97.5 31.8 ;
      RECT 91.5 30.6 97.5 31.8 ;
      RECT 87.9 28.2 89.1 29.4 ;
      RECT 87.9 5.1 88.8 29.4 ;
      RECT 87.6 15.9 88.8 17.1 ;
      RECT 87.9 5.1 89.1 6.3 ;
      RECT 85.2 29.1 86.4 31.8 ;
      RECT 85.5 13.8 86.4 31.8 ;
      RECT 85.2 18.3 86.4 19.5 ;
      RECT 85.2 13.8 86.4 15 ;
      RECT 82.2 31.5 83.4 33.3 ;
      RECT 82.5 11.7 83.4 33.3 ;
      RECT 82.5 26.7 83.7 27.9 ;
      RECT 82.2 20.7 83.4 21.9 ;
      RECT 82.5 11.7 83.7 12.9 ;
      RECT 79.2 33.9 80.4 35.7 ;
      RECT 79.2 9.6 80.1 35.7 ;
      RECT 79.2 23.1 80.4 24.3 ;
      RECT 79.2 9.6 80.4 10.8 ;
      RECT 76.8 28.2 78 29.4 ;
      RECT 77.1 5.1 78 29.4 ;
      RECT 76.8 15.9 78 17.1 ;
      RECT 77.1 5.1 78.3 6.3 ;
      RECT 71.1 6.6 74.1 7.8 ;
      RECT 75 6 76.2 7.2 ;
      RECT 73.2 6.3 76.2 7.2 ;
      RECT 71.1 14.4 74.1 15.9 ;
      RECT 71.1 14.4 75.3 15.3 ;
      RECT 75.3 8.1 76.2 14.7 ;
      RECT 74.1 13.8 76.2 14.7 ;
      RECT 75 8.1 76.2 9.3 ;
      RECT 71.1 21.9 74.1 23.1 ;
      RECT 71.1 21.9 75.9 22.8 ;
      RECT 75 17.4 75.9 22.8 ;
      RECT 71.1 17.4 75.9 18.3 ;
      RECT 71.1 17.1 74.1 18.3 ;
      RECT 71.1 35.4 74.1 36.6 ;
      RECT 71.1 35.4 75.9 36.3 ;
      RECT 75 30.9 75.9 36.3 ;
      RECT 71.1 30.9 75.9 31.8 ;
      RECT 71.1 30.6 74.1 31.8 ;
      RECT 64.2 0.6 70.2 36.9 ;
      RECT 60.3 33 74.1 34.2 ;
      RECT 60.3 24.3 74.1 25.5 ;
      RECT 60.3 19.5 74.1 20.7 ;
      RECT 60.3 9 74.1 10.2 ;
      RECT 60.3 4.2 74.1 5.4 ;
      RECT 60.3 6.6 63.3 7.8 ;
      RECT 58.2 6.3 61.2 7.2 ;
      RECT 58.2 6 59.4 7.2 ;
      RECT 60.3 14.4 63.3 15.9 ;
      RECT 59.1 13.8 60.3 15.3 ;
      RECT 58.2 8.1 59.1 14.7 ;
      RECT 58.2 8.1 59.4 9.3 ;
      RECT 60.3 21.9 63.3 23.1 ;
      RECT 58.5 21.9 63.3 22.8 ;
      RECT 58.5 17.4 59.4 22.8 ;
      RECT 58.5 17.4 63.3 18.3 ;
      RECT 60.3 17.1 63.3 18.3 ;
      RECT 60.3 35.4 63.3 36.6 ;
      RECT 58.5 35.4 63.3 36.3 ;
      RECT 58.5 30.9 59.4 36.3 ;
      RECT 58.5 30.9 63.3 31.8 ;
      RECT 60.3 30.6 63.3 31.8 ;
      RECT 56.4 28.2 57.6 29.4 ;
      RECT 56.4 5.1 57.3 29.4 ;
      RECT 56.4 15.9 57.6 17.1 ;
      RECT 56.1 5.1 57.3 6.3 ;
      RECT 54 33.9 55.2 35.7 ;
      RECT 54.3 9.6 55.2 35.7 ;
      RECT 54 23.1 55.2 24.3 ;
      RECT 54 9.6 55.2 10.8 ;
      RECT 51 31.5 52.2 33.3 ;
      RECT 51 11.7 51.9 33.3 ;
      RECT 50.7 26.7 51.9 27.9 ;
      RECT 51 20.7 52.2 21.9 ;
      RECT 50.7 11.7 51.9 12.9 ;
      RECT 48 29.1 49.2 31.8 ;
      RECT 48 13.8 48.9 31.8 ;
      RECT 48 18.3 49.2 19.5 ;
      RECT 48 13.8 49.2 15 ;
      RECT 45.3 28.2 46.5 29.4 ;
      RECT 45.6 5.1 46.5 29.4 ;
      RECT 45.6 15.9 46.8 17.1 ;
      RECT 45.3 5.1 46.5 6.3 ;
      RECT 36.9 21.9 42.9 23.1 ;
      RECT 36.9 21.9 44.7 22.8 ;
      RECT 43.8 17.4 44.7 22.8 ;
      RECT 36.9 17.4 44.7 18.3 ;
      RECT 36.9 17.1 42.9 18.3 ;
      RECT 36.9 35.4 42.9 36.6 ;
      RECT 36.9 35.4 44.7 36.3 ;
      RECT 43.8 30.9 44.7 36.3 ;
      RECT 36.9 30.9 44.7 31.8 ;
      RECT 36.9 30.6 42.9 31.8 ;
      RECT 36.9 14.4 42.9 15.9 ;
      RECT 42 13.8 44.1 15 ;
      RECT 35.1 0.6 36 37.2 ;
      RECT 35.1 33 42.9 34.2 ;
      RECT 35.1 24.3 42.9 25.5 ;
      RECT 35.1 19.5 42.9 20.7 ;
      RECT 35.1 9 42.9 10.2 ;
      RECT 35.1 4.2 42.9 5.4 ;
      RECT 31.2 0.6 32.1 37.2 ;
      RECT 24.3 33 32.1 34.2 ;
      RECT 24.3 24.3 32.1 25.5 ;
      RECT 24.3 19.5 32.1 20.7 ;
      RECT 24.3 9 32.1 10.2 ;
      RECT 24.3 4.2 32.1 5.4 ;
      RECT 24.3 14.4 30.3 15.9 ;
      RECT 23.1 13.8 25.2 15 ;
      RECT 24.3 21.9 30.3 23.1 ;
      RECT 22.5 21.9 30.3 22.8 ;
      RECT 22.5 17.4 23.4 22.8 ;
      RECT 22.5 17.4 30.3 18.3 ;
      RECT 24.3 17.1 30.3 18.3 ;
      RECT 24.3 35.4 30.3 36.6 ;
      RECT 22.5 35.4 30.3 36.3 ;
      RECT 22.5 30.9 23.4 36.3 ;
      RECT 22.5 30.9 30.3 31.8 ;
      RECT 24.3 30.6 30.3 31.8 ;
      RECT 20.7 28.2 21.9 29.4 ;
      RECT 20.7 5.1 21.6 29.4 ;
      RECT 20.4 15.9 21.6 17.1 ;
      RECT 20.7 5.1 21.9 6.3 ;
      RECT 18 29.1 19.2 30.9 ;
      RECT 18.3 13.8 19.2 30.9 ;
      RECT 18 18.3 19.2 19.5 ;
      RECT 18 13.8 19.2 15 ;
      RECT 15 31.5 16.2 33.3 ;
      RECT 15.3 11.7 16.2 33.3 ;
      RECT 15.3 26.7 16.5 27.9 ;
      RECT 15 20.7 16.2 21.9 ;
      RECT 15.3 11.7 16.5 12.9 ;
      RECT 12 33.9 13.2 35.7 ;
      RECT 12 9.6 12.9 35.7 ;
      RECT 12 23.1 13.2 24.3 ;
      RECT 12 9.6 13.2 10.8 ;
      RECT 9.6 28.2 10.8 29.4 ;
      RECT 9.9 5.1 10.8 29.4 ;
      RECT 9.6 15.9 10.8 17.1 ;
      RECT 9.9 5.1 11.1 6.3 ;
      RECT 3.9 6.6 6.9 7.8 ;
      RECT 7.8 6 9 7.2 ;
      RECT 6 6.3 9 7.2 ;
      RECT 3.9 14.4 6.9 15.9 ;
      RECT 3.9 14.4 8.1 15.3 ;
      RECT 8.1 8.1 9 14.7 ;
      RECT 6.9 13.8 9 14.7 ;
      RECT 7.8 8.1 9 9.3 ;
      RECT 3.9 21.9 6.9 23.1 ;
      RECT 3.9 21.9 8.7 22.8 ;
      RECT 7.8 17.4 8.7 22.8 ;
      RECT 3.9 17.4 8.7 18.3 ;
      RECT 3.9 17.1 6.9 18.3 ;
      RECT 3.9 35.4 6.9 36.6 ;
      RECT 3.9 35.4 8.7 36.3 ;
      RECT 7.8 30.9 8.7 36.3 ;
      RECT 3.9 30.9 8.7 31.8 ;
      RECT 3.9 30.6 6.9 31.8 ;
      RECT 260.7 1.8 264.9 3 ;
      RECT 261.9 4.2 264.9 5.4 ;
      RECT 261.9 9 264.9 10.2 ;
      RECT 261.9 19.5 264.9 20.7 ;
      RECT 261.9 24.3 264.9 25.5 ;
      RECT 260.7 28.2 264.9 29.4 ;
      RECT 261.9 33 264.9 34.2 ;
      RECT 255.6 2.7 256.8 3 ;
      RECT 252.6 1.5 253.8 7.8 ;
      RECT 238.5 1.8 245.7 3 ;
      RECT 238.5 6.6 245.7 7.8 ;
      RECT 238.5 28.2 245.7 29.4 ;
      RECT 224.7 1.8 231.9 3 ;
      RECT 224.7 6.6 231.9 7.8 ;
      RECT 224.7 28.2 231.9 29.4 ;
      RECT 216.6 1.5 217.8 7.8 ;
      RECT 213.6 1.8 214.8 3 ;
      RECT 205.5 1.8 209.7 3 ;
      RECT 205.5 28.2 209.7 29.4 ;
      RECT 193.5 1.8 197.7 3 ;
      RECT 193.5 28.2 197.7 29.4 ;
      RECT 188.4 1.8 189.6 3 ;
      RECT 185.4 1.5 186.6 7.8 ;
      RECT 171.3 1.8 178.5 3 ;
      RECT 171.3 6.6 178.5 7.8 ;
      RECT 171.3 28.2 178.5 29.4 ;
      RECT 157.5 1.8 164.7 3 ;
      RECT 157.5 6.6 164.7 7.8 ;
      RECT 157.5 28.2 164.7 29.4 ;
      RECT 149.4 1.5 150.6 7.8 ;
      RECT 146.4 1.8 147.6 3 ;
      RECT 138.3 1.8 142.5 3 ;
      RECT 138.3 28.2 142.5 29.4 ;
      RECT 126.3 1.8 130.5 3 ;
      RECT 126.3 28.2 130.5 29.4 ;
      RECT 121.2 1.8 122.4 3 ;
      RECT 118.2 1.5 119.4 7.8 ;
      RECT 104.1 1.8 111.3 3 ;
      RECT 104.1 6.6 111.3 7.8 ;
      RECT 104.1 28.2 111.3 29.4 ;
      RECT 90.3 1.8 97.5 3 ;
      RECT 90.3 6.6 97.5 7.8 ;
      RECT 90.3 28.2 97.5 29.4 ;
      RECT 82.2 1.5 83.4 7.8 ;
      RECT 79.2 1.8 80.4 3 ;
      RECT 71.1 1.8 75.3 3 ;
      RECT 71.1 28.2 75.3 29.4 ;
      RECT 59.1 1.8 63.3 3 ;
      RECT 59.1 28.2 63.3 29.4 ;
      RECT 54 1.8 55.2 3 ;
      RECT 51 1.5 52.2 7.8 ;
      RECT 36.9 1.8 44.1 3 ;
      RECT 36.9 6.6 44.1 7.8 ;
      RECT 36.9 28.2 44.1 29.4 ;
      RECT 23.1 1.8 30.3 3 ;
      RECT 23.1 6.6 30.3 7.8 ;
      RECT 23.1 28.2 30.3 29.4 ;
      RECT 15 1.5 16.2 7.8 ;
      RECT 12 1.8 13.2 3 ;
      RECT 3.9 1.8 8.1 3 ;
      RECT 3.9 28.2 8.1 29.4 ;
      RECT 3.9 4.2 6.9 5.4 ;
      RECT 3.9 9 6.9 10.2 ;
      RECT 3.9 19.5 6.9 20.7 ;
      RECT 3.9 24.3 6.9 25.5 ;
      RECT 3.9 33 6.9 34.2 ;
  END
END rca8

END LIBRARY
