/home/dshadoa/Desktop/BPM/chip/abstract/bpm_custom.lef