* SPICE NETLIST
***************************************

.SUBCKT dffpos clk_b D clk Q
** N=21 EP=4 IP=0 FDC=26
M0 16 clk_b 8 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=9900 $Y=19500 $D=1
M1 clk clk_b 16 8 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=11400 $Y=19500 $D=1
M2 17 D 8 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=16200 $Y=19500 $D=1
M3 4 clk_b 17 8 n L=6e-07 W=3e-06 AD=5.4e-12 AS=2.7e-12 PD=9.6e-06 PS=7.8e-06 $X=17700 $Y=19500 $D=1
M4 18 clk 4 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=5.4e-12 PD=7.8e-06 PS=9.6e-06 $X=20100 $Y=19500 $D=1
M5 8 5 18 8 n L=6e-07 W=3e-06 AD=6.3e-12 AS=2.7e-12 PD=1.02e-05 PS=7.8e-06 $X=21600 $Y=19500 $D=1
M6 5 4 8 8 n L=6e-07 W=3e-06 AD=4.5e-12 AS=6.3e-12 PD=9e-06 PS=1.02e-05 $X=24300 $Y=19500 $D=1
M7 19 5 8 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=29100 $Y=19500 $D=1
M8 6 clk 19 8 n L=6e-07 W=3e-06 AD=5.4e-12 AS=2.7e-12 PD=9.6e-06 PS=7.8e-06 $X=30600 $Y=19500 $D=1
M9 20 clk_b 6 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=5.4e-12 PD=7.8e-06 PS=9.6e-06 $X=33000 $Y=19500 $D=1
M10 8 Q 20 8 n L=6e-07 W=3e-06 AD=6.3e-12 AS=2.7e-12 PD=1.02e-05 PS=7.8e-06 $X=34500 $Y=19500 $D=1
M11 21 6 8 8 n L=6e-07 W=3e-06 AD=2.7e-12 AS=6.3e-12 PD=7.8e-06 PS=1.02e-05 $X=37200 $Y=19500 $D=1
M12 Q 6 21 8 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=38700 $Y=19500 $D=1
M13 10 clk_b 7 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=9900 $Y=2700 $D=0
M14 clk clk_b 10 7 p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=11400 $Y=2700 $D=0
M15 11 D 7 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=16200 $Y=2700 $D=0
M16 4 clk 11 7 p L=6e-07 W=6e-06 AD=1.08e-11 AS=5.4e-12 PD=1.56e-05 PS=1.38e-05 $X=17700 $Y=2700 $D=0
M17 12 clk_b 4 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.08e-11 PD=1.38e-05 PS=1.56e-05 $X=20100 $Y=2700 $D=0
M18 7 5 12 7 p L=6e-07 W=6e-06 AD=1.26e-11 AS=5.4e-12 PD=1.62e-05 PS=1.38e-05 $X=21600 $Y=2700 $D=0
M19 5 4 7 7 p L=6e-07 W=6e-06 AD=9e-12 AS=1.26e-11 PD=1.5e-05 PS=1.62e-05 $X=24300 $Y=2700 $D=0
M20 13 5 7 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=29100 $Y=2700 $D=0
M21 6 clk_b 13 7 p L=6e-07 W=6e-06 AD=1.08e-11 AS=5.4e-12 PD=1.56e-05 PS=1.38e-05 $X=30600 $Y=2700 $D=0
M22 14 clk 6 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.08e-11 PD=1.38e-05 PS=1.56e-05 $X=33000 $Y=2700 $D=0
M23 7 Q 14 7 p L=6e-07 W=6e-06 AD=1.26e-11 AS=5.4e-12 PD=1.62e-05 PS=1.38e-05 $X=34500 $Y=2700 $D=0
M24 15 6 7 7 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.26e-11 PD=1.38e-05 PS=1.62e-05 $X=37200 $Y=2700 $D=0
M25 Q 6 15 7 p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=38700 $Y=2700 $D=0
.ENDS
***************************************
