magic
tech scmos
timestamp 1542302220
<< ntransistor >>
rect 96 65 98 75
<< ptransistor >>
rect 96 9 98 29
<< ndiffusion >>
rect 95 65 96 75
rect 98 65 99 75
<< pdiffusion >>
rect 95 9 96 29
rect 98 9 99 29
<< ndcontact >>
rect 91 65 95 75
rect 99 65 103 75
<< pdcontact >>
rect 91 9 95 29
rect 99 9 103 29
<< psubstratepcontact >>
rect 87 79 91 83
rect 103 79 107 83
<< nsubstratencontact >>
rect 88 1 92 5
rect 102 1 106 5
<< polysilicon >>
rect 96 75 98 77
rect 96 58 98 65
rect 95 54 98 58
rect 96 29 98 54
rect 96 7 98 9
<< polycontact >>
rect 91 54 95 58
<< metal1 >>
rect -1 174 244 177
rect 64 168 69 174
rect 236 168 244 174
rect -1 145 8 149
rect 64 83 244 96
rect 64 79 87 83
rect 91 79 103 83
rect 107 79 244 83
rect 64 78 244 79
rect 91 75 95 78
rect 86 54 91 58
rect 73 48 74 52
rect 99 29 103 65
rect -1 24 8 28
rect -1 17 8 21
rect 91 6 95 9
rect -1 5 244 6
rect -1 1 88 5
rect 92 1 102 5
rect 106 1 244 5
rect -1 -3 244 1
<< m2contact >>
rect 8 145 12 149
rect 74 48 78 52
rect 67 38 71 42
rect 8 24 12 28
rect 8 17 12 21
<< metal2 >>
rect 12 145 79 149
rect 75 123 79 145
rect 75 119 88 123
rect 60 112 67 116
rect 60 102 64 112
rect 64 71 108 75
rect 67 28 71 38
rect 12 24 71 28
rect 74 21 78 48
rect 12 17 78 21
use ../../fa/magic/fa  fa_0 ../../fa/magic
timestamp 1542251572
transform 1 0 61 0 1 90
box 0 -4 175 89
use ../../bc1a/magic/bc1a  bc1a_0 ../../bc1a/magic
timestamp 1542169151
transform 1 0 0 0 1 12
box -1 -12 64 162
use ../../nand/magic/nand  nand_0 ../../nand/magic
timestamp 1542301814
transform 1 0 65 0 -1 81
box -4 -3 28 81
<< labels >>
rlabel metal1 176 176 176 176 5 c_in
rlabel metal1 1 147 1 147 3 fa_in
rlabel metal1 1 26 1 26 3 clk
rlabel metal1 1 19 1 19 3 en
rlabel metal2 106 73 106 73 1 from_mux
rlabel metal1 101 48 101 48 1 from_and
<< end >>
