magic
tech scmos
timestamp 1542725905
<< metal1 >>
rect -4 2 0 129
rect 36 122 40 129
rect 46 114 50 129
rect 106 2 110 129
rect 166 114 170 129
rect 176 122 180 129
rect 216 2 220 129
<< metal2 >>
rect 94 103 156 106
rect 94 9 97 103
rect 77 6 97 9
use fa  fa_0
timestamp 1541616290
transform 0 1 3 -1 0 124
box -5 -3 124 105
use fa  fa_1
timestamp 1541616290
transform 0 -1 213 -1 0 124
box -5 -3 124 105
<< end >>
