magic
tech scmos
timestamp 1542725905
<< metal1 >>
rect -3 2 3 3
rect -3 -2 -2 2
rect 2 -2 3 2
rect -3 -3 3 -2
<< m2contact >>
rect -2 -2 2 2
<< metal2 >>
rect -3 2 3 3
rect -3 -2 -2 2
rect 2 -2 3 2
rect -3 -3 3 -2
<< end >>
