magic
tech scmos
timestamp 1543290821
<< ntransistor >>
rect 11 9 13 19
rect 19 9 21 19
rect 35 9 37 19
rect 51 9 53 19
rect 56 9 58 19
rect 72 9 74 19
rect 80 9 82 19
rect 88 9 90 19
rect 104 9 106 19
rect 120 9 122 19
rect 125 9 127 19
rect 130 9 132 19
rect 146 9 148 19
rect 162 9 164 19
<< ptransistor >>
rect 11 55 13 75
rect 19 55 21 75
rect 35 55 37 75
rect 51 55 53 75
rect 56 55 58 75
rect 72 55 74 75
rect 80 55 82 75
rect 88 55 90 75
rect 104 55 106 75
rect 120 55 122 75
rect 125 55 127 75
rect 130 55 132 75
rect 146 55 148 75
rect 162 55 164 75
<< ndiffusion >>
rect 10 9 11 19
rect 13 9 14 19
rect 18 9 19 19
rect 21 9 22 19
rect 34 9 35 19
rect 37 9 38 19
rect 50 9 51 19
rect 53 9 56 19
rect 58 9 59 19
rect 71 9 72 19
rect 74 9 75 19
rect 79 9 80 19
rect 82 9 83 19
rect 87 9 88 19
rect 90 9 91 19
rect 103 9 104 19
rect 106 9 107 19
rect 119 9 120 19
rect 122 9 125 19
rect 127 9 130 19
rect 132 9 133 19
rect 145 9 146 19
rect 148 9 149 19
rect 161 9 162 19
rect 164 9 165 19
<< pdiffusion >>
rect 10 55 11 75
rect 13 55 14 75
rect 18 55 19 75
rect 21 55 22 75
rect 34 55 35 75
rect 37 55 38 75
rect 50 55 51 75
rect 53 55 56 75
rect 58 55 59 75
rect 71 55 72 75
rect 74 55 75 75
rect 79 55 80 75
rect 82 55 83 75
rect 87 55 88 75
rect 90 55 91 75
rect 103 55 104 75
rect 106 55 107 75
rect 119 55 120 75
rect 122 55 125 75
rect 127 55 130 75
rect 132 55 133 75
rect 145 55 146 75
rect 148 55 149 75
rect 161 55 162 75
rect 164 55 165 75
<< ndcontact >>
rect 6 9 10 19
rect 14 9 18 19
rect 22 9 26 19
rect 30 9 34 19
rect 38 9 42 19
rect 46 9 50 19
rect 59 9 63 19
rect 67 9 71 19
rect 75 9 79 19
rect 83 9 87 19
rect 91 9 95 19
rect 99 9 103 19
rect 107 9 111 19
rect 115 9 119 19
rect 133 9 137 19
rect 141 9 145 19
rect 149 9 153 19
rect 157 9 161 19
rect 165 9 169 19
<< pdcontact >>
rect 6 55 10 75
rect 14 55 18 75
rect 22 55 26 75
rect 30 55 34 75
rect 38 55 42 75
rect 46 55 50 75
rect 59 55 63 75
rect 67 55 71 75
rect 75 55 79 75
rect 83 55 87 75
rect 91 55 95 75
rect 99 55 103 75
rect 107 55 111 75
rect 115 55 119 75
rect 133 55 137 75
rect 141 55 145 75
rect 149 55 153 75
rect 157 55 161 75
rect 165 55 169 75
<< psubstratepcontact >>
rect 10 1 14 5
rect 18 1 22 5
rect 34 1 38 5
rect 46 1 50 5
rect 59 1 63 5
rect 71 1 75 5
rect 79 1 83 5
rect 87 1 91 5
rect 103 1 107 5
rect 115 1 119 5
rect 124 1 128 5
rect 133 1 137 5
rect 149 1 153 5
rect 165 1 169 5
<< nsubstratencontact >>
rect 10 79 14 83
rect 18 79 22 83
rect 34 79 38 83
rect 46 79 50 83
rect 59 79 63 83
rect 71 79 75 83
rect 79 79 83 83
rect 87 79 91 83
rect 103 79 107 83
rect 115 79 119 83
rect 124 79 128 83
rect 133 79 137 83
rect 149 79 153 83
rect 165 79 169 83
<< polysilicon >>
rect 11 75 13 77
rect 19 75 21 77
rect 35 75 37 77
rect 51 75 53 77
rect 56 75 58 77
rect 72 75 74 77
rect 80 75 82 77
rect 88 75 90 77
rect 104 75 106 77
rect 120 75 122 77
rect 125 75 127 77
rect 130 75 132 77
rect 146 75 148 77
rect 162 75 164 77
rect 11 30 13 55
rect 10 26 13 30
rect 11 19 13 26
rect 19 33 21 55
rect 35 45 37 55
rect 34 41 37 45
rect 51 44 53 55
rect 19 29 22 33
rect 19 19 21 29
rect 35 19 37 41
rect 50 40 53 44
rect 51 36 53 40
rect 46 34 53 36
rect 46 22 48 34
rect 46 20 53 22
rect 51 19 53 20
rect 56 19 58 55
rect 72 52 74 55
rect 71 48 74 52
rect 72 19 74 48
rect 80 48 82 55
rect 88 54 90 55
rect 88 52 95 54
rect 80 46 85 48
rect 83 33 85 46
rect 82 29 85 33
rect 83 24 85 29
rect 80 22 85 24
rect 93 22 95 52
rect 104 40 106 55
rect 120 54 122 55
rect 103 36 106 40
rect 80 19 82 22
rect 88 20 95 22
rect 88 19 90 20
rect 104 19 106 36
rect 115 52 122 54
rect 115 22 117 52
rect 120 40 121 44
rect 125 40 127 55
rect 120 27 122 40
rect 120 25 127 27
rect 115 20 122 22
rect 120 19 122 20
rect 125 19 127 25
rect 130 19 132 55
rect 146 26 148 55
rect 162 33 164 55
rect 161 29 164 33
rect 145 22 148 26
rect 146 19 148 22
rect 162 19 164 29
rect 11 7 13 9
rect 19 7 21 9
rect 35 7 37 9
rect 51 7 53 9
rect 56 7 58 9
rect 72 7 74 9
rect 80 7 82 9
rect 88 7 90 9
rect 104 7 106 9
rect 120 7 122 9
rect 125 7 127 9
rect 130 7 132 9
rect 146 7 148 9
rect 162 7 164 9
<< polycontact >>
rect 6 26 10 30
rect 30 41 34 45
rect 22 29 26 33
rect 46 40 50 44
rect 52 26 56 30
rect 67 48 71 52
rect 78 29 82 33
rect 89 29 93 33
rect 99 36 103 40
rect 117 48 121 52
rect 121 40 125 44
rect 126 32 130 36
rect 157 29 161 33
rect 141 22 145 26
<< metal1 >>
rect 0 83 175 84
rect 0 79 10 83
rect 14 79 18 83
rect 22 79 34 83
rect 38 79 46 83
rect 50 79 59 83
rect 63 79 71 83
rect 75 79 79 83
rect 83 79 87 83
rect 91 79 103 83
rect 107 79 115 83
rect 119 79 124 83
rect 128 79 133 83
rect 137 79 149 83
rect 153 79 165 83
rect 169 79 175 83
rect 0 78 175 79
rect 6 75 10 78
rect 22 75 26 78
rect 46 75 50 78
rect 67 75 71 78
rect 83 75 87 78
rect 115 75 119 78
rect 141 75 145 78
rect 157 75 161 78
rect 14 52 18 55
rect 30 52 34 55
rect 14 48 34 52
rect 38 52 42 55
rect 59 52 63 55
rect 75 52 79 55
rect 91 52 95 55
rect 99 52 103 55
rect 38 48 63 52
rect 14 22 34 26
rect 14 19 18 22
rect 30 19 34 22
rect 38 19 42 48
rect 59 40 63 48
rect 75 48 103 52
rect 59 36 99 40
rect 59 19 63 36
rect 99 33 103 36
rect 71 29 78 33
rect 107 29 110 55
rect 134 29 137 55
rect 107 26 137 29
rect 149 52 153 55
rect 75 22 103 26
rect 75 19 79 22
rect 91 19 95 22
rect 99 19 103 22
rect 107 19 110 26
rect 134 22 141 26
rect 134 19 137 22
rect 149 19 153 48
rect 165 19 169 55
rect 6 6 10 9
rect 22 6 26 9
rect 46 6 50 9
rect 67 6 71 9
rect 83 6 87 9
rect 115 6 119 9
rect 141 6 145 9
rect 157 6 161 9
rect 0 5 175 6
rect 0 1 10 5
rect 14 1 18 5
rect 22 1 34 5
rect 38 1 46 5
rect 50 1 59 5
rect 63 1 71 5
rect 75 1 79 5
rect 83 1 87 5
rect 91 1 103 5
rect 107 1 115 5
rect 119 1 124 5
rect 128 1 133 5
rect 137 1 149 5
rect 153 1 165 5
rect 169 1 175 5
rect 0 0 175 1
<< m2contact >>
rect 26 41 30 45
rect 26 29 30 33
rect 6 22 10 26
rect 46 36 50 40
rect 67 44 71 48
rect 52 22 56 26
rect 67 29 71 33
rect 85 29 89 33
rect 99 29 103 33
rect 113 48 117 52
rect 117 40 121 44
rect 122 32 126 36
rect 149 48 153 52
rect 157 25 161 29
rect 169 22 173 26
<< metal2 >>
rect 113 55 117 87
rect 67 52 117 55
rect 67 51 113 52
rect 67 48 71 51
rect 153 48 175 52
rect 26 45 67 48
rect 30 44 67 45
rect 74 45 110 48
rect 74 44 121 45
rect 74 40 78 44
rect 107 42 117 44
rect 39 36 46 40
rect 50 36 78 40
rect 85 36 114 39
rect 39 33 43 36
rect 30 29 43 33
rect 67 33 71 36
rect 85 33 89 36
rect 85 26 89 29
rect 10 22 52 26
rect 56 22 89 26
rect 111 32 122 36
rect 99 25 157 29
rect 169 -4 173 22
<< labels >>
rlabel metal1 3 81 3 81 4 vdd
rlabel metal1 3 3 3 3 3 gnd
rlabel polysilicon 12 39 12 39 1 a
rlabel polysilicon 20 39 20 39 1 b
rlabel metal2 112 53 112 53 5 c_in
rlabel metal2 159 50 159 50 7 sum
rlabel metal2 171 20 171 20 8 c_out
<< end >>
