/classes/ecen4303F18/osu_soc_3.0/lib/ami05/lib/osu05_stdcells.lef