magic
tech scmos
timestamp 1543295583
<< ntransistor >>
rect 36 43 38 53
rect 44 43 46 53
<< ptransistor >>
rect 36 7 38 17
rect 44 7 46 17
<< ndiffusion >>
rect 35 43 36 53
rect 38 43 39 53
rect 43 43 44 53
rect 46 43 47 53
<< pdiffusion >>
rect 35 7 36 17
rect 38 7 39 17
rect 43 7 44 17
rect 46 7 47 17
<< ndcontact >>
rect 31 43 35 53
rect 39 43 43 53
rect 47 43 51 53
<< pdcontact >>
rect 31 7 35 17
rect 39 7 43 17
rect 47 7 51 17
<< psubstratepcontact >>
rect 39 67 43 71
rect 49 67 53 71
<< nsubstratencontact >>
rect 31 -11 35 -7
rect 48 -11 52 -7
<< polysilicon >>
rect 36 58 54 60
rect 36 53 38 58
rect 44 53 46 55
rect 36 41 38 43
rect 44 38 46 43
rect 36 36 46 38
rect 36 17 38 36
rect 44 18 54 20
rect 44 17 46 18
rect 36 2 38 7
rect 44 5 46 7
<< polycontact >>
rect 54 57 58 61
rect 54 17 58 21
rect 36 -2 40 2
<< metal1 >>
rect -1 156 30 162
rect 46 156 61 162
rect -1 148 1 152
rect 5 148 20 152
rect 23 118 27 122
rect 38 93 42 97
rect -1 87 12 91
rect -1 83 30 84
rect -1 79 28 83
rect 42 80 61 84
rect -1 78 30 79
rect 33 78 64 80
rect -1 72 64 78
rect -1 71 58 72
rect -1 66 9 71
rect 30 67 39 71
rect 43 67 49 71
rect 53 67 58 71
rect 30 66 58 67
rect 39 53 43 59
rect -1 37 8 41
rect 31 34 35 43
rect -1 30 8 34
rect 23 26 27 30
rect 31 17 35 30
rect 39 17 43 43
rect 47 41 51 43
rect 47 17 51 37
rect 54 50 58 57
rect 54 21 58 46
rect -1 -12 9 -6
rect 30 -7 58 -6
rect 30 -11 31 -7
rect 35 -11 48 -7
rect 52 -11 64 -7
rect 30 -12 64 -11
<< m2contact >>
rect 1 148 5 152
rect 38 87 42 91
rect 39 59 43 63
rect 8 46 12 50
rect 23 46 27 50
rect 8 37 12 41
rect 8 30 12 34
rect 31 30 35 34
rect 47 37 51 41
rect 54 46 58 50
rect 32 -2 36 2
<< metal2 >>
rect 1 50 5 148
rect 38 77 42 87
rect 32 73 42 77
rect 32 50 36 73
rect 43 59 58 63
rect 1 46 8 50
rect 27 46 54 50
rect 1 2 5 46
rect 12 37 47 41
rect 12 30 31 34
rect 30 12 62 16
rect 30 5 62 9
rect 1 -2 32 2
use mux21  mux21_0
timestamp 1543295496
transform 1 0 38 0 1 115
box -30 -37 4 47
use inverter  inverter_1
timestamp 1543289418
transform 1 0 13 0 -1 71
box -4 -1 20 83
<< labels >>
rlabel metal2 14 32 14 32 3 a_in
rlabel metal2 14 39 14 39 3 b_in
rlabel metal1 8 75 8 75 3 gnd
rlabel metal1 7 89 7 89 3 reg_in
<< end >>
