magic
tech scmos
timestamp 1542725905
<< m2contact >>
rect -2 -2 2 2
<< end >>
