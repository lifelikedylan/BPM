magic
tech scmos
timestamp 1543282798
<< metal1 >>
rect -1 174 218 177
rect 61 168 218 174
rect -1 145 4 149
rect 58 89 218 96
rect 64 83 218 89
rect 64 78 87 83
rect 93 78 218 83
rect 86 54 87 58
rect 73 48 74 52
rect 199 42 218 47
rect -1 24 8 28
rect -1 17 8 21
rect -1 1 87 6
rect 93 1 218 6
rect -1 -3 218 1
<< m2contact >>
rect 4 145 8 149
rect 74 48 78 52
rect 67 38 71 42
rect 8 24 12 28
rect 8 17 12 21
<< metal2 >>
rect 8 145 48 149
rect 201 82 216 86
rect 201 81 206 82
rect 64 71 87 75
rect 67 28 71 38
rect 12 24 71 28
rect 74 21 78 48
rect 12 17 78 21
rect 201 4 205 81
rect 156 0 205 4
rect 156 -3 160 0
use ../../bc1a/magic/bc1a  bc1a_0 ../../bc1a/magic
timestamp 1543282357
transform 1 0 0 0 1 12
box -1 -12 64 162
use ../../nand/magic/nand  nand_0 ../../nand/magic
timestamp 1543271335
transform 1 0 65 0 -1 81
box -4 -3 28 81
use ../../dffpos/magic/dffpos  dffpos_0 ../../dffpos/magic
timestamp 1543271063
transform 1 0 63 0 1 0
box 18 0 139 84
<< labels >>
rlabel metal1 1 26 1 26 3 clk
rlabel metal1 1 19 1 19 3 en
rlabel metal1 5 1 5 1 1 vdd
rlabel space 5 173 5 173 5 vdd
rlabel metal1 1 147 1 147 3 fa_in
rlabel space 1 114 1 114 3 Init
rlabel space 0 101 0 101 3 reg_in
rlabel metal1 216 45 216 45 7 Out
rlabel space 0 51 0 51 3 muxB_in
rlabel space 0 44 0 44 3 muxA_in
rlabel space -2 86 -2 86 3 gnd
rlabel metal1 158 -2 158 -2 1 Cout
<< end >>
