magic
tech scmos
magscale 1 2
timestamp 1542725905
<< metal1 >>
rect -10 4 10 6
rect -10 -4 -9 4
rect 9 -4 10 4
rect -10 -6 10 -4
<< m2contact >>
rect -9 -4 9 4
<< metal2 >>
rect -10 4 10 6
rect -10 -4 -9 4
rect 9 -4 10 4
rect -10 -6 10 -4
<< end >>
