VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO bpm_custom
  CLASS RING ;
  ORIGIN 4.8 18.3 ;
  FOREIGN bpm_custom -4.8 -18.3 ;
  SIZE 162.6 BY 457.2 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 -5.4 82.2 -3.6 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 -2.7 80.1 -0.9 ;
    END
  END en
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER metal2 ;
        RECT 52.8 432.9 77.7 434.1 ;
      LAYER metal1 ;
        RECT 26.4 25.8 86.4 29.7 ;
        RECT 35.1 24.3 86.4 29.7 ;
        RECT 26.4 24.3 33.3 29.7 ;
        RECT 26.4 403.8 86.4 407.7 ;
        RECT 35.1 402.3 86.4 407.7 ;
        RECT 26.4 402.3 33.3 407.7 ;
        RECT 0 -8.1 78 -6.3 ;
    END
  END gnd
  PIN init
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 -13.5 88.5 -11.7 ;
    END
  END init
  PIN mcand_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 417.3 153 418.5 ;
    END
  END mcand_0
  PIN mcand_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 363.3 153 364.5 ;
    END
  END mcand_1
  PIN mcand_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 309.3 153 310.5 ;
    END
  END mcand_2
  PIN mcand_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 255.3 153 256.5 ;
    END
  END mcand_3
  PIN mcand_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 201.3 153 202.5 ;
    END
  END mcand_4
  PIN mcand_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 147.3 153 148.5 ;
    END
  END mcand_5
  PIN mcand_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 93.3 153 94.5 ;
    END
  END mcand_6
  PIN mcand_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 39.3 153 40.5 ;
    END
  END mcand_7
  PIN mplier_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 415.2 153 416.4 ;
    END
  END mplier_0
  PIN mplier_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 361.2 153 362.4 ;
    END
  END mplier_1
  PIN mplier_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 307.2 153 308.4 ;
    END
  END mplier_2
  PIN mplier_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 253.2 153 254.4 ;
    END
  END mplier_3
  PIN mplier_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 199.2 153 200.4 ;
    END
  END mplier_4
  PIN mplier_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 145.2 153 146.4 ;
    END
  END mplier_5
  PIN mplier_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 91.2 153 92.4 ;
    END
  END mplier_6
  PIN mplier_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114 37.2 153 38.4 ;
    END
  END mplier_7
  PIN q_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 391.5 153 393 ;
    END
  END q_0
  PIN q_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 337.5 153 339 ;
    END
  END q_1
  PIN q_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 288.3 72.9 289.5 ;
    END
  END q_10
  PIN q_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 234.3 72.9 235.5 ;
    END
  END q_11
  PIN q_12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 180.3 72.9 181.5 ;
    END
  END q_12
  PIN q_13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 126.3 72.9 127.5 ;
    END
  END q_13
  PIN q_14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 72.3 72.9 73.5 ;
    END
  END q_14
  PIN q_15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 18.3 72.9 19.5 ;
    END
  END q_15
  PIN q_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 283.5 153 285 ;
    END
  END q_2
  PIN q_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 229.5 153 231 ;
    END
  END q_3
  PIN q_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 175.5 153 177 ;
    END
  END q_4
  PIN q_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 121.5 153 123 ;
    END
  END q_5
  PIN q_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 67.5 153 69 ;
    END
  END q_6
  PIN q_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 144.6 13.5 153 15 ;
    END
  END q_7
  PIN q_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 396.3 72.9 397.5 ;
    END
  END q_8
  PIN q_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.9 342.3 72.9 343.5 ;
    END
  END q_9
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER metal1 ;
        RECT 114.6 0 153 2.7 ;
        RECT 0 0 153 1.2 ;
        RECT 35.1 0 112.8 2.7 ;
        RECT 0 0 33.3 2.7 ;
        RECT 0 431.1 153 432 ;
        RECT 99 429.3 153 432 ;
        RECT 71.1 429.3 86.4 432 ;
        RECT 26.4 429.3 27.9 432 ;
        RECT 0 429.3 6.9 432 ;
        RECT 0 -10.8 75.9 -9 ;
        RECT 26.4 51.3 27.9 56.7 ;
        RECT 26.4 105.3 27.9 110.7 ;
        RECT 26.4 159.3 27.9 164.7 ;
        RECT 26.4 213.3 27.9 218.7 ;
        RECT 26.4 267.3 27.9 272.7 ;
        RECT 26.4 321.3 27.9 326.7 ;
        RECT 26.4 375.3 27.9 380.7 ;
    END
  END vdd
  PIN cout
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.8 0 54 0.9 ;
    END
  END cout
  OBS
    LAYER metal2 ;
      RECT 91.2 34.5 150.9 35.7 ;
      RECT 149.7 13.5 150.9 35.7 ;
      RECT 91.2 30.6 92.4 35.7 ;
      RECT 91.2 88.5 150.9 89.7 ;
      RECT 149.7 67.5 150.9 89.7 ;
      RECT 91.2 84.6 92.4 89.7 ;
      RECT 91.2 142.5 150.9 143.7 ;
      RECT 149.7 121.5 150.9 143.7 ;
      RECT 91.2 138.6 92.4 143.7 ;
      RECT 91.2 196.5 150.9 197.7 ;
      RECT 149.7 175.5 150.9 197.7 ;
      RECT 91.2 192.6 92.4 197.7 ;
      RECT 91.2 250.5 150.9 251.7 ;
      RECT 149.7 229.5 150.9 251.7 ;
      RECT 91.2 246.6 92.4 251.7 ;
      RECT 91.2 304.5 150.9 305.7 ;
      RECT 149.7 283.5 150.9 305.7 ;
      RECT 91.2 300.6 92.4 305.7 ;
      RECT 91.2 358.5 150.9 359.7 ;
      RECT 149.7 337.5 150.9 359.7 ;
      RECT 91.2 354.6 92.4 359.7 ;
      RECT 91.2 412.5 150.9 413.7 ;
      RECT 149.7 391.5 150.9 413.7 ;
      RECT 91.2 408.6 92.4 413.7 ;
      RECT 131.7 15.9 137.1 17.1 ;
      RECT 135.9 10.5 137.1 17.1 ;
      RECT 120.6 10.5 137.1 11.7 ;
      RECT 131.7 69.9 137.1 71.1 ;
      RECT 135.9 64.5 137.1 71.1 ;
      RECT 120.6 64.5 137.1 65.7 ;
      RECT 131.7 123.9 137.1 125.1 ;
      RECT 135.9 118.5 137.1 125.1 ;
      RECT 120.6 118.5 137.1 119.7 ;
      RECT 131.7 177.9 137.1 179.1 ;
      RECT 135.9 172.5 137.1 179.1 ;
      RECT 120.6 172.5 137.1 173.7 ;
      RECT 131.7 231.9 137.1 233.1 ;
      RECT 135.9 226.5 137.1 233.1 ;
      RECT 120.6 226.5 137.1 227.7 ;
      RECT 131.7 285.9 137.1 287.1 ;
      RECT 135.9 280.5 137.1 287.1 ;
      RECT 120.6 280.5 137.1 281.7 ;
      RECT 131.7 339.9 137.1 341.1 ;
      RECT 135.9 334.5 137.1 341.1 ;
      RECT 120.6 334.5 137.1 335.7 ;
      RECT 131.7 393.9 137.1 395.1 ;
      RECT 135.9 388.5 137.1 395.1 ;
      RECT 120.6 388.5 137.1 389.7 ;
      RECT 113.7 18.3 121.8 19.5 ;
      RECT 120.6 14.4 121.8 19.5 ;
      RECT 120.6 14.4 130.2 15.6 ;
      RECT 129 13.5 133.5 14.7 ;
      RECT 113.7 72.3 121.8 73.5 ;
      RECT 120.6 68.4 121.8 73.5 ;
      RECT 120.6 68.4 130.2 69.6 ;
      RECT 129 67.5 133.5 68.7 ;
      RECT 113.7 126.3 121.8 127.5 ;
      RECT 120.6 122.4 121.8 127.5 ;
      RECT 120.6 122.4 130.2 123.6 ;
      RECT 129 121.5 133.5 122.7 ;
      RECT 113.7 180.3 121.8 181.5 ;
      RECT 120.6 176.4 121.8 181.5 ;
      RECT 120.6 176.4 130.2 177.6 ;
      RECT 129 175.5 133.5 176.7 ;
      RECT 113.7 234.3 121.8 235.5 ;
      RECT 120.6 230.4 121.8 235.5 ;
      RECT 120.6 230.4 130.2 231.6 ;
      RECT 129 229.5 133.5 230.7 ;
      RECT 113.7 288.3 121.8 289.5 ;
      RECT 120.6 284.4 121.8 289.5 ;
      RECT 120.6 284.4 130.2 285.6 ;
      RECT 129 283.5 133.5 284.7 ;
      RECT 113.7 342.3 121.8 343.5 ;
      RECT 120.6 338.4 121.8 343.5 ;
      RECT 120.6 338.4 130.2 339.6 ;
      RECT 129 337.5 133.5 338.7 ;
      RECT 113.7 396.3 121.8 397.5 ;
      RECT 120.6 392.4 121.8 397.5 ;
      RECT 120.6 392.4 130.2 393.6 ;
      RECT 129 391.5 133.5 392.7 ;
      RECT 98.4 22.2 112.8 23.4 ;
      RECT 111.6 14.7 112.8 23.4 ;
      RECT 111.6 14.7 119.4 15.9 ;
      RECT 98.4 76.2 112.8 77.4 ;
      RECT 111.6 68.7 112.8 77.4 ;
      RECT 111.6 68.7 119.4 69.9 ;
      RECT 98.4 130.2 112.8 131.4 ;
      RECT 111.6 122.7 112.8 131.4 ;
      RECT 111.6 122.7 119.4 123.9 ;
      RECT 98.4 184.2 112.8 185.4 ;
      RECT 111.6 176.7 112.8 185.4 ;
      RECT 111.6 176.7 119.4 177.9 ;
      RECT 98.4 238.2 112.8 239.4 ;
      RECT 111.6 230.7 112.8 239.4 ;
      RECT 111.6 230.7 119.4 231.9 ;
      RECT 98.4 292.2 112.8 293.4 ;
      RECT 111.6 284.7 112.8 293.4 ;
      RECT 111.6 284.7 119.4 285.9 ;
      RECT 98.4 346.2 112.8 347.4 ;
      RECT 111.6 338.7 112.8 347.4 ;
      RECT 111.6 338.7 119.4 339.9 ;
      RECT 98.4 400.2 112.8 401.4 ;
      RECT 111.6 392.7 112.8 401.4 ;
      RECT 111.6 392.7 119.4 393.9 ;
      RECT 107.4 29.7 108.6 33.6 ;
      RECT 107.4 29.7 108.9 31.2 ;
      RECT 107.4 83.7 108.6 87.6 ;
      RECT 107.4 83.7 108.9 85.2 ;
      RECT 107.4 137.7 108.6 141.6 ;
      RECT 107.4 137.7 108.9 139.2 ;
      RECT 107.4 191.7 108.6 195.6 ;
      RECT 107.4 191.7 108.9 193.2 ;
      RECT 107.4 245.7 108.6 249.6 ;
      RECT 107.4 245.7 108.9 247.2 ;
      RECT 107.4 299.7 108.6 303.6 ;
      RECT 107.4 299.7 108.9 301.2 ;
      RECT 107.4 353.7 108.6 357.6 ;
      RECT 107.4 353.7 108.9 355.2 ;
      RECT 107.4 407.7 108.6 411.6 ;
      RECT 107.4 407.7 108.9 409.2 ;
      RECT 107.1 6 108.3 16.5 ;
      RECT 89.1 6 108.3 7.2 ;
      RECT 107.1 60 108.3 70.5 ;
      RECT 89.1 60 108.3 61.2 ;
      RECT 107.1 114 108.3 124.5 ;
      RECT 89.1 114 108.3 115.2 ;
      RECT 107.1 168 108.3 178.5 ;
      RECT 89.1 168 108.3 169.2 ;
      RECT 107.1 222 108.3 232.5 ;
      RECT 89.1 222 108.3 223.2 ;
      RECT 107.1 276 108.3 286.5 ;
      RECT 89.1 276 108.3 277.2 ;
      RECT 107.1 330 108.3 340.5 ;
      RECT 89.1 330 108.3 331.2 ;
      RECT 107.1 384 108.3 394.5 ;
      RECT 89.1 384 108.3 385.2 ;
      RECT 100.5 48.9 106.5 50.1 ;
      RECT 100.5 41.4 101.7 50.1 ;
      RECT 89.1 41.4 101.7 42.6 ;
      RECT 100.5 102.9 106.5 104.1 ;
      RECT 100.5 95.4 101.7 104.1 ;
      RECT 89.1 95.4 101.7 96.6 ;
      RECT 100.5 156.9 106.5 158.1 ;
      RECT 100.5 149.4 101.7 158.1 ;
      RECT 89.1 149.4 101.7 150.6 ;
      RECT 100.5 210.9 106.5 212.1 ;
      RECT 100.5 203.4 101.7 212.1 ;
      RECT 89.1 203.4 101.7 204.6 ;
      RECT 100.5 264.9 106.5 266.1 ;
      RECT 100.5 257.4 101.7 266.1 ;
      RECT 89.1 257.4 101.7 258.6 ;
      RECT 100.5 318.9 106.5 320.1 ;
      RECT 100.5 311.4 101.7 320.1 ;
      RECT 89.1 311.4 101.7 312.6 ;
      RECT 100.5 372.9 106.5 374.1 ;
      RECT 100.5 365.4 101.7 374.1 ;
      RECT 89.1 365.4 101.7 366.6 ;
      RECT 100.5 426.9 106.5 428.1 ;
      RECT 100.5 419.4 101.7 428.1 ;
      RECT 89.1 419.4 101.7 420.6 ;
      RECT 105 8.1 106.2 13.5 ;
      RECT 89.1 8.1 106.2 9.3 ;
      RECT 105 62.1 106.2 67.5 ;
      RECT 89.1 62.1 106.2 63.3 ;
      RECT 105 116.1 106.2 121.5 ;
      RECT 89.1 116.1 106.2 117.3 ;
      RECT 105 170.1 106.2 175.5 ;
      RECT 89.1 170.1 106.2 171.3 ;
      RECT 105 224.1 106.2 229.5 ;
      RECT 89.1 224.1 106.2 225.3 ;
      RECT 105 278.1 106.2 283.5 ;
      RECT 89.1 278.1 106.2 279.3 ;
      RECT 105 332.1 106.2 337.5 ;
      RECT 89.1 332.1 106.2 333.3 ;
      RECT 105 386.1 106.2 391.5 ;
      RECT 89.1 386.1 106.2 387.3 ;
      RECT 98.1 26.4 99.3 31.8 ;
      RECT 96.3 26.4 99.3 27.6 ;
      RECT 96.3 18.3 97.5 27.6 ;
      RECT 93.6 18.3 104.1 19.5 ;
      RECT 98.1 80.4 99.3 85.8 ;
      RECT 96.3 80.4 99.3 81.6 ;
      RECT 96.3 72.3 97.5 81.6 ;
      RECT 93.6 72.3 104.1 73.5 ;
      RECT 98.1 134.4 99.3 139.8 ;
      RECT 96.3 134.4 99.3 135.6 ;
      RECT 96.3 126.3 97.5 135.6 ;
      RECT 93.6 126.3 104.1 127.5 ;
      RECT 98.1 188.4 99.3 193.8 ;
      RECT 96.3 188.4 99.3 189.6 ;
      RECT 96.3 180.3 97.5 189.6 ;
      RECT 93.6 180.3 104.1 181.5 ;
      RECT 98.1 242.4 99.3 247.8 ;
      RECT 96.3 242.4 99.3 243.6 ;
      RECT 96.3 234.3 97.5 243.6 ;
      RECT 93.6 234.3 104.1 235.5 ;
      RECT 98.1 296.4 99.3 301.8 ;
      RECT 96.3 296.4 99.3 297.6 ;
      RECT 96.3 288.3 97.5 297.6 ;
      RECT 93.6 288.3 104.1 289.5 ;
      RECT 98.1 350.4 99.3 355.8 ;
      RECT 96.3 350.4 99.3 351.6 ;
      RECT 96.3 342.3 97.5 351.6 ;
      RECT 93.6 342.3 104.1 343.5 ;
      RECT 98.1 404.4 99.3 409.8 ;
      RECT 96.3 404.4 99.3 405.6 ;
      RECT 96.3 396.3 97.5 405.6 ;
      RECT 93.6 396.3 104.1 397.5 ;
      RECT 93.6 26.4 94.8 33.6 ;
      RECT 91.2 26.4 94.8 27.6 ;
      RECT 91.2 15.6 92.4 27.6 ;
      RECT 89.1 15.6 102 16.8 ;
      RECT 93.6 80.4 94.8 87.6 ;
      RECT 91.2 80.4 94.8 81.6 ;
      RECT 91.2 69.6 92.4 81.6 ;
      RECT 89.1 69.6 102 70.8 ;
      RECT 93.6 134.4 94.8 141.6 ;
      RECT 91.2 134.4 94.8 135.6 ;
      RECT 91.2 123.6 92.4 135.6 ;
      RECT 89.1 123.6 102 124.8 ;
      RECT 93.6 188.4 94.8 195.6 ;
      RECT 91.2 188.4 94.8 189.6 ;
      RECT 91.2 177.6 92.4 189.6 ;
      RECT 89.1 177.6 102 178.8 ;
      RECT 93.6 242.4 94.8 249.6 ;
      RECT 91.2 242.4 94.8 243.6 ;
      RECT 91.2 231.6 92.4 243.6 ;
      RECT 89.1 231.6 102 232.8 ;
      RECT 93.6 296.4 94.8 303.6 ;
      RECT 91.2 296.4 94.8 297.6 ;
      RECT 91.2 285.6 92.4 297.6 ;
      RECT 89.1 285.6 102 286.8 ;
      RECT 93.6 350.4 94.8 357.6 ;
      RECT 91.2 350.4 94.8 351.6 ;
      RECT 91.2 339.6 92.4 351.6 ;
      RECT 89.1 339.6 102 340.8 ;
      RECT 93.6 404.4 94.8 411.6 ;
      RECT 91.2 404.4 94.8 405.6 ;
      RECT 91.2 393.6 92.4 405.6 ;
      RECT 89.1 393.6 102 394.8 ;
      RECT 87 -13.2 88.2 432 ;
      RECT 87 396.3 90.3 397.5 ;
      RECT 87 381.9 97.5 383.1 ;
      RECT 87 342.3 90.3 343.5 ;
      RECT 87 327.9 97.5 329.1 ;
      RECT 87 288.3 90.3 289.5 ;
      RECT 87 273.9 97.5 275.1 ;
      RECT 87 234.3 90.3 235.5 ;
      RECT 87 219.9 97.5 221.1 ;
      RECT 87 180.3 90.3 181.5 ;
      RECT 87 165.9 97.5 167.1 ;
      RECT 87 126.3 90.3 127.5 ;
      RECT 87 111.9 97.5 113.1 ;
      RECT 87 72.3 90.3 73.5 ;
      RECT 87 57.9 97.5 59.1 ;
      RECT 87 18.3 90.3 19.5 ;
      RECT 87 3.9 97.5 5.1 ;
      RECT 84.9 -2.4 86.1 14.7 ;
      RECT 84.6 -2.4 86.1 -0.9 ;
      RECT 41.1 41.1 51.9 42.3 ;
      RECT 41.1 41.1 55.2 41.4 ;
      RECT 71.1 39.6 72.6 41.1 ;
      RECT 54 39.9 72.6 41.1 ;
      RECT 51 40.5 72.6 41.1 ;
      RECT 41.1 38.7 42.3 42.3 ;
      RECT 30.6 38.7 42.3 39.9 ;
      RECT 39 36.6 40.2 39.9 ;
      RECT 30.6 36.6 31.8 39.9 ;
      RECT 26.7 36.6 31.8 37.8 ;
      RECT 41.1 95.1 51.9 96.3 ;
      RECT 41.1 95.1 55.2 95.4 ;
      RECT 71.1 93.6 72.6 95.1 ;
      RECT 54 93.9 72.6 95.1 ;
      RECT 51 94.5 72.6 95.1 ;
      RECT 41.1 92.7 42.3 96.3 ;
      RECT 30.6 92.7 42.3 93.9 ;
      RECT 39 90.6 40.2 93.9 ;
      RECT 30.6 90.6 31.8 93.9 ;
      RECT 26.7 90.6 31.8 91.8 ;
      RECT 41.1 149.1 51.9 150.3 ;
      RECT 41.1 149.1 55.2 149.4 ;
      RECT 71.1 147.6 72.6 149.1 ;
      RECT 54 147.9 72.6 149.1 ;
      RECT 51 148.5 72.6 149.1 ;
      RECT 41.1 146.7 42.3 150.3 ;
      RECT 30.6 146.7 42.3 147.9 ;
      RECT 39 144.6 40.2 147.9 ;
      RECT 30.6 144.6 31.8 147.9 ;
      RECT 26.7 144.6 31.8 145.8 ;
      RECT 41.1 203.1 51.9 204.3 ;
      RECT 41.1 203.1 55.2 203.4 ;
      RECT 71.1 201.6 72.6 203.1 ;
      RECT 54 201.9 72.6 203.1 ;
      RECT 51 202.5 72.6 203.1 ;
      RECT 41.1 200.7 42.3 204.3 ;
      RECT 30.6 200.7 42.3 201.9 ;
      RECT 39 198.6 40.2 201.9 ;
      RECT 30.6 198.6 31.8 201.9 ;
      RECT 26.7 198.6 31.8 199.8 ;
      RECT 41.1 257.1 51.9 258.3 ;
      RECT 41.1 257.1 55.2 257.4 ;
      RECT 71.1 255.6 72.6 257.1 ;
      RECT 54 255.9 72.6 257.1 ;
      RECT 51 256.5 72.6 257.1 ;
      RECT 41.1 254.7 42.3 258.3 ;
      RECT 30.6 254.7 42.3 255.9 ;
      RECT 39 252.6 40.2 255.9 ;
      RECT 30.6 252.6 31.8 255.9 ;
      RECT 26.7 252.6 31.8 253.8 ;
      RECT 41.1 311.1 51.9 312.3 ;
      RECT 41.1 311.1 55.2 311.4 ;
      RECT 71.1 309.6 72.6 311.1 ;
      RECT 54 309.9 72.6 311.1 ;
      RECT 51 310.5 72.6 311.1 ;
      RECT 41.1 308.7 42.3 312.3 ;
      RECT 30.6 308.7 42.3 309.9 ;
      RECT 39 306.6 40.2 309.9 ;
      RECT 30.6 306.6 31.8 309.9 ;
      RECT 26.7 306.6 31.8 307.8 ;
      RECT 41.1 365.1 51.9 366.3 ;
      RECT 41.1 365.1 55.2 365.4 ;
      RECT 71.1 363.6 72.6 365.1 ;
      RECT 54 363.9 72.6 365.1 ;
      RECT 51 364.5 72.6 365.1 ;
      RECT 41.1 362.7 42.3 366.3 ;
      RECT 30.6 362.7 42.3 363.9 ;
      RECT 39 360.6 40.2 363.9 ;
      RECT 30.6 360.6 31.8 363.9 ;
      RECT 26.7 360.6 31.8 361.8 ;
      RECT 41.1 419.1 51.9 420.3 ;
      RECT 41.1 419.1 55.2 419.4 ;
      RECT 71.1 417.6 72.6 419.1 ;
      RECT 54 417.9 72.6 419.1 ;
      RECT 51 418.5 72.6 419.1 ;
      RECT 41.1 416.7 42.3 420.3 ;
      RECT 30.6 416.7 42.3 417.9 ;
      RECT 39 414.6 40.2 417.9 ;
      RECT 30.6 414.6 31.8 417.9 ;
      RECT 26.7 414.6 31.8 415.8 ;
      RECT 68.1 52.2 69.6 53.7 ;
      RECT 68.4 42.3 69.6 53.7 ;
      RECT 63.6 42.3 71.4 43.5 ;
      RECT 68.1 106.2 69.6 107.7 ;
      RECT 68.4 96.3 69.6 107.7 ;
      RECT 63.6 96.3 71.4 97.5 ;
      RECT 68.1 160.2 69.6 161.7 ;
      RECT 68.4 150.3 69.6 161.7 ;
      RECT 63.6 150.3 71.4 151.5 ;
      RECT 68.1 214.2 69.6 215.7 ;
      RECT 68.4 204.3 69.6 215.7 ;
      RECT 63.6 204.3 71.4 205.5 ;
      RECT 68.1 268.2 69.6 269.7 ;
      RECT 68.4 258.3 69.6 269.7 ;
      RECT 63.6 258.3 71.4 259.5 ;
      RECT 68.1 322.2 69.6 323.7 ;
      RECT 68.4 312.3 69.6 323.7 ;
      RECT 63.6 312.3 71.4 313.5 ;
      RECT 68.1 376.2 69.6 377.7 ;
      RECT 68.4 366.3 69.6 377.7 ;
      RECT 63.6 366.3 71.4 367.5 ;
      RECT 68.1 430.2 69.6 431.7 ;
      RECT 68.4 420.3 69.6 431.7 ;
      RECT 63.6 420.3 71.4 421.5 ;
      RECT 69.6 0.9 70.8 35.7 ;
      RECT 68.1 0.9 70.8 3.6 ;
      RECT 52.8 1.8 70.8 2.1 ;
      RECT 54.9 0.9 70.8 2.1 ;
      RECT 69.6 54.9 70.8 89.7 ;
      RECT 52.8 54.9 70.8 56.1 ;
      RECT 52.8 42.3 54 56.1 ;
      RECT 39 43.2 54 44.4 ;
      RECT 39 41.1 40.2 44.4 ;
      RECT 26.7 41.1 40.2 42.3 ;
      RECT 26.7 40.2 27.9 42.3 ;
      RECT 69.6 108.9 70.8 143.7 ;
      RECT 52.8 108.9 70.8 110.1 ;
      RECT 52.8 96.3 54 110.1 ;
      RECT 39 97.2 54 98.4 ;
      RECT 39 95.1 40.2 98.4 ;
      RECT 26.7 95.1 40.2 96.3 ;
      RECT 26.7 94.2 27.9 96.3 ;
      RECT 69.6 162.9 70.8 197.7 ;
      RECT 52.8 162.9 70.8 164.1 ;
      RECT 52.8 150.3 54 164.1 ;
      RECT 39 151.2 54 152.4 ;
      RECT 39 149.1 40.2 152.4 ;
      RECT 26.7 149.1 40.2 150.3 ;
      RECT 26.7 148.2 27.9 150.3 ;
      RECT 69.6 216.9 70.8 251.7 ;
      RECT 52.8 216.9 70.8 218.1 ;
      RECT 52.8 204.3 54 218.1 ;
      RECT 39 205.2 54 206.4 ;
      RECT 39 203.1 40.2 206.4 ;
      RECT 26.7 203.1 40.2 204.3 ;
      RECT 26.7 202.2 27.9 204.3 ;
      RECT 69.6 270.9 70.8 305.7 ;
      RECT 52.8 270.9 70.8 272.1 ;
      RECT 52.8 258.3 54 272.1 ;
      RECT 39 259.2 54 260.4 ;
      RECT 39 257.1 40.2 260.4 ;
      RECT 26.7 257.1 40.2 258.3 ;
      RECT 26.7 256.2 27.9 258.3 ;
      RECT 69.6 324.9 70.8 359.7 ;
      RECT 52.8 324.9 70.8 326.1 ;
      RECT 52.8 312.3 54 326.1 ;
      RECT 39 313.2 54 314.4 ;
      RECT 39 311.1 40.2 314.4 ;
      RECT 26.7 311.1 40.2 312.3 ;
      RECT 26.7 310.2 27.9 312.3 ;
      RECT 69.6 378.9 70.8 413.7 ;
      RECT 52.8 378.9 70.8 380.1 ;
      RECT 52.8 366.3 54 380.1 ;
      RECT 39 367.2 54 368.4 ;
      RECT 39 365.1 40.2 368.4 ;
      RECT 26.7 365.1 40.2 366.3 ;
      RECT 26.7 364.2 27.9 366.3 ;
      RECT 48.6 35.4 49.8 37.8 ;
      RECT 48.6 35.4 67.2 36.6 ;
      RECT 48.6 89.4 49.8 91.8 ;
      RECT 48.6 89.4 67.2 90.6 ;
      RECT 48.6 143.4 49.8 145.8 ;
      RECT 48.6 143.4 67.2 144.6 ;
      RECT 48.6 197.4 49.8 199.8 ;
      RECT 48.6 197.4 67.2 198.6 ;
      RECT 48.6 251.4 49.8 253.8 ;
      RECT 48.6 251.4 67.2 252.6 ;
      RECT 48.6 305.4 49.8 307.8 ;
      RECT 48.6 305.4 67.2 306.6 ;
      RECT 48.6 359.4 49.8 361.8 ;
      RECT 48.6 359.4 67.2 360.6 ;
      RECT 48.6 413.4 49.8 415.8 ;
      RECT 48.6 413.4 67.2 414.6 ;
      RECT 11.7 32.7 21.9 33.6 ;
      RECT 20.7 26.4 21.9 33.6 ;
      RECT 11.7 32.4 17.7 33.6 ;
      RECT 20.7 26.4 65.1 27.6 ;
      RECT 63.9 18.3 65.1 27.6 ;
      RECT 11.7 86.7 21.9 87.6 ;
      RECT 20.7 80.4 21.9 87.6 ;
      RECT 11.7 86.4 17.7 87.6 ;
      RECT 20.7 80.4 65.1 81.6 ;
      RECT 63.9 72.3 65.1 81.6 ;
      RECT 11.7 140.7 21.9 141.6 ;
      RECT 20.7 134.4 21.9 141.6 ;
      RECT 11.7 140.4 17.7 141.6 ;
      RECT 20.7 134.4 65.1 135.6 ;
      RECT 63.9 126.3 65.1 135.6 ;
      RECT 11.7 194.7 21.9 195.6 ;
      RECT 20.7 188.4 21.9 195.6 ;
      RECT 11.7 194.4 17.7 195.6 ;
      RECT 20.7 188.4 65.1 189.6 ;
      RECT 63.9 180.3 65.1 189.6 ;
      RECT 11.7 248.7 21.9 249.6 ;
      RECT 20.7 242.4 21.9 249.6 ;
      RECT 11.7 248.4 17.7 249.6 ;
      RECT 20.7 242.4 65.1 243.6 ;
      RECT 63.9 234.3 65.1 243.6 ;
      RECT 11.7 302.7 21.9 303.6 ;
      RECT 20.7 296.4 21.9 303.6 ;
      RECT 11.7 302.4 17.7 303.6 ;
      RECT 20.7 296.4 65.1 297.6 ;
      RECT 63.9 288.3 65.1 297.6 ;
      RECT 11.7 356.7 21.9 357.6 ;
      RECT 20.7 350.4 21.9 357.6 ;
      RECT 11.7 356.4 17.7 357.6 ;
      RECT 20.7 350.4 65.1 351.6 ;
      RECT 63.9 342.3 65.1 351.6 ;
      RECT 11.7 410.7 21.9 411.6 ;
      RECT 20.7 404.4 21.9 411.6 ;
      RECT 11.7 410.4 17.7 411.6 ;
      RECT 20.7 404.4 65.1 405.6 ;
      RECT 63.9 396.3 65.1 405.6 ;
      RECT 52.2 15.9 57.6 17.1 ;
      RECT 56.4 10.5 57.6 17.1 ;
      RECT 41.1 10.5 57.6 11.7 ;
      RECT 52.2 69.9 57.6 71.1 ;
      RECT 56.4 64.5 57.6 71.1 ;
      RECT 41.1 64.5 57.6 65.7 ;
      RECT 52.2 123.9 57.6 125.1 ;
      RECT 56.4 118.5 57.6 125.1 ;
      RECT 41.1 118.5 57.6 119.7 ;
      RECT 52.2 177.9 57.6 179.1 ;
      RECT 56.4 172.5 57.6 179.1 ;
      RECT 41.1 172.5 57.6 173.7 ;
      RECT 52.2 231.9 57.6 233.1 ;
      RECT 56.4 226.5 57.6 233.1 ;
      RECT 41.1 226.5 57.6 227.7 ;
      RECT 52.2 285.9 57.6 287.1 ;
      RECT 56.4 280.5 57.6 287.1 ;
      RECT 41.1 280.5 57.6 281.7 ;
      RECT 52.2 339.9 57.6 341.1 ;
      RECT 56.4 334.5 57.6 341.1 ;
      RECT 41.1 334.5 57.6 335.7 ;
      RECT 52.2 393.9 57.6 395.1 ;
      RECT 56.4 388.5 57.6 395.1 ;
      RECT 41.1 388.5 57.6 389.7 ;
      RECT 14.1 39.3 21.9 40.5 ;
      RECT 20.7 34.5 21.9 40.5 ;
      RECT 44.4 38.7 53.1 39.6 ;
      RECT 52.2 37.5 56.7 38.7 ;
      RECT 44.4 34.5 45.6 39.6 ;
      RECT 20.7 34.5 45.6 35.7 ;
      RECT 14.1 93.3 21.9 94.5 ;
      RECT 20.7 88.5 21.9 94.5 ;
      RECT 44.4 92.7 53.1 93.6 ;
      RECT 52.2 91.5 56.7 92.7 ;
      RECT 44.4 88.5 45.6 93.6 ;
      RECT 20.7 88.5 45.6 89.7 ;
      RECT 14.1 147.3 21.9 148.5 ;
      RECT 20.7 142.5 21.9 148.5 ;
      RECT 44.4 146.7 53.1 147.6 ;
      RECT 52.2 145.5 56.7 146.7 ;
      RECT 44.4 142.5 45.6 147.6 ;
      RECT 20.7 142.5 45.6 143.7 ;
      RECT 14.1 201.3 21.9 202.5 ;
      RECT 20.7 196.5 21.9 202.5 ;
      RECT 44.4 200.7 53.1 201.6 ;
      RECT 52.2 199.5 56.7 200.7 ;
      RECT 44.4 196.5 45.6 201.6 ;
      RECT 20.7 196.5 45.6 197.7 ;
      RECT 14.1 255.3 21.9 256.5 ;
      RECT 20.7 250.5 21.9 256.5 ;
      RECT 44.4 254.7 53.1 255.6 ;
      RECT 52.2 253.5 56.7 254.7 ;
      RECT 44.4 250.5 45.6 255.6 ;
      RECT 20.7 250.5 45.6 251.7 ;
      RECT 14.1 309.3 21.9 310.5 ;
      RECT 20.7 304.5 21.9 310.5 ;
      RECT 44.4 308.7 53.1 309.6 ;
      RECT 52.2 307.5 56.7 308.7 ;
      RECT 44.4 304.5 45.6 309.6 ;
      RECT 20.7 304.5 45.6 305.7 ;
      RECT 14.1 363.3 21.9 364.5 ;
      RECT 20.7 358.5 21.9 364.5 ;
      RECT 44.4 362.7 53.1 363.6 ;
      RECT 52.2 361.5 56.7 362.7 ;
      RECT 44.4 358.5 45.6 363.6 ;
      RECT 20.7 358.5 45.6 359.7 ;
      RECT 14.1 417.3 21.9 418.5 ;
      RECT 20.7 412.5 21.9 418.5 ;
      RECT 44.4 416.7 53.1 417.6 ;
      RECT 52.2 415.5 56.7 416.7 ;
      RECT 44.4 412.5 45.6 417.6 ;
      RECT 20.7 412.5 45.6 413.7 ;
      RECT 34.2 18.3 42.3 19.5 ;
      RECT 41.1 14.4 42.3 19.5 ;
      RECT 41.1 14.4 50.7 15.6 ;
      RECT 49.5 13.5 54 14.7 ;
      RECT 34.2 72.3 42.3 73.5 ;
      RECT 41.1 68.4 42.3 73.5 ;
      RECT 41.1 68.4 50.7 69.6 ;
      RECT 49.5 67.5 54 68.7 ;
      RECT 34.2 126.3 42.3 127.5 ;
      RECT 41.1 122.4 42.3 127.5 ;
      RECT 41.1 122.4 50.7 123.6 ;
      RECT 49.5 121.5 54 122.7 ;
      RECT 34.2 180.3 42.3 181.5 ;
      RECT 41.1 176.4 42.3 181.5 ;
      RECT 41.1 176.4 50.7 177.6 ;
      RECT 49.5 175.5 54 176.7 ;
      RECT 34.2 234.3 42.3 235.5 ;
      RECT 41.1 230.4 42.3 235.5 ;
      RECT 41.1 230.4 50.7 231.6 ;
      RECT 49.5 229.5 54 230.7 ;
      RECT 34.2 288.3 42.3 289.5 ;
      RECT 41.1 284.4 42.3 289.5 ;
      RECT 41.1 284.4 50.7 285.6 ;
      RECT 49.5 283.5 54 284.7 ;
      RECT 34.2 342.3 42.3 343.5 ;
      RECT 41.1 338.4 42.3 343.5 ;
      RECT 41.1 338.4 50.7 339.6 ;
      RECT 49.5 337.5 54 338.7 ;
      RECT 34.2 396.3 42.3 397.5 ;
      RECT 41.1 392.4 42.3 397.5 ;
      RECT 41.1 392.4 50.7 393.6 ;
      RECT 49.5 391.5 54 392.7 ;
      RECT 52.8 420.3 54 432 ;
      RECT 39 421.2 54 422.4 ;
      RECT 39 419.1 40.2 422.4 ;
      RECT 26.7 419.1 40.2 420.3 ;
      RECT 26.7 418.2 27.9 420.3 ;
      RECT 18.9 22.2 33.3 23.4 ;
      RECT 32.1 14.7 33.3 23.4 ;
      RECT 32.1 14.7 39.9 15.9 ;
      RECT 18.9 76.2 33.3 77.4 ;
      RECT 32.1 68.7 33.3 77.4 ;
      RECT 32.1 68.7 39.9 69.9 ;
      RECT 18.9 130.2 33.3 131.4 ;
      RECT 32.1 122.7 33.3 131.4 ;
      RECT 32.1 122.7 39.9 123.9 ;
      RECT 18.9 184.2 33.3 185.4 ;
      RECT 32.1 176.7 33.3 185.4 ;
      RECT 32.1 176.7 39.9 177.9 ;
      RECT 18.9 238.2 33.3 239.4 ;
      RECT 32.1 230.7 33.3 239.4 ;
      RECT 32.1 230.7 39.9 231.9 ;
      RECT 18.9 292.2 33.3 293.4 ;
      RECT 32.1 284.7 33.3 293.4 ;
      RECT 32.1 284.7 39.9 285.9 ;
      RECT 18.9 346.2 33.3 347.4 ;
      RECT 32.1 338.7 33.3 347.4 ;
      RECT 32.1 338.7 39.9 339.9 ;
      RECT 18.9 400.2 33.3 401.4 ;
      RECT 32.1 392.7 33.3 401.4 ;
      RECT 32.1 392.7 39.9 393.9 ;
      RECT 27.6 6 28.8 16.5 ;
      RECT 9.6 6 28.8 7.2 ;
      RECT 27.6 60 28.8 70.5 ;
      RECT 9.6 60 28.8 61.2 ;
      RECT 27.6 114 28.8 124.5 ;
      RECT 9.6 114 28.8 115.2 ;
      RECT 27.6 168 28.8 178.5 ;
      RECT 9.6 168 28.8 169.2 ;
      RECT 27.6 222 28.8 232.5 ;
      RECT 9.6 222 28.8 223.2 ;
      RECT 27.6 276 28.8 286.5 ;
      RECT 9.6 276 28.8 277.2 ;
      RECT 27.6 330 28.8 340.5 ;
      RECT 9.6 330 28.8 331.2 ;
      RECT 27.6 384 28.8 394.5 ;
      RECT 9.6 384 28.8 385.2 ;
      RECT 25.5 8.1 26.7 13.5 ;
      RECT 9.6 8.1 26.7 9.3 ;
      RECT 25.5 62.1 26.7 67.5 ;
      RECT 9.6 62.1 26.7 63.3 ;
      RECT 25.5 116.1 26.7 121.5 ;
      RECT 9.6 116.1 26.7 117.3 ;
      RECT 25.5 170.1 26.7 175.5 ;
      RECT 9.6 170.1 26.7 171.3 ;
      RECT 25.5 224.1 26.7 229.5 ;
      RECT 9.6 224.1 26.7 225.3 ;
      RECT 25.5 278.1 26.7 283.5 ;
      RECT 9.6 278.1 26.7 279.3 ;
      RECT 25.5 332.1 26.7 337.5 ;
      RECT 9.6 332.1 26.7 333.3 ;
      RECT 25.5 386.1 26.7 391.5 ;
      RECT 9.6 386.1 26.7 387.3 ;
      RECT 18.6 26.4 19.8 31.8 ;
      RECT 16.8 26.4 19.8 27.6 ;
      RECT 16.8 18.3 18 27.6 ;
      RECT 14.1 18.3 24.6 19.5 ;
      RECT 18.6 80.4 19.8 85.8 ;
      RECT 16.8 80.4 19.8 81.6 ;
      RECT 16.8 72.3 18 81.6 ;
      RECT 14.1 72.3 24.6 73.5 ;
      RECT 18.6 134.4 19.8 139.8 ;
      RECT 16.8 134.4 19.8 135.6 ;
      RECT 16.8 126.3 18 135.6 ;
      RECT 14.1 126.3 24.6 127.5 ;
      RECT 18.6 188.4 19.8 193.8 ;
      RECT 16.8 188.4 19.8 189.6 ;
      RECT 16.8 180.3 18 189.6 ;
      RECT 14.1 180.3 24.6 181.5 ;
      RECT 18.6 242.4 19.8 247.8 ;
      RECT 16.8 242.4 19.8 243.6 ;
      RECT 16.8 234.3 18 243.6 ;
      RECT 14.1 234.3 24.6 235.5 ;
      RECT 18.6 296.4 19.8 301.8 ;
      RECT 16.8 296.4 19.8 297.6 ;
      RECT 16.8 288.3 18 297.6 ;
      RECT 14.1 288.3 24.6 289.5 ;
      RECT 18.6 350.4 19.8 355.8 ;
      RECT 16.8 350.4 19.8 351.6 ;
      RECT 16.8 342.3 18 351.6 ;
      RECT 14.1 342.3 24.6 343.5 ;
      RECT 18.6 404.4 19.8 409.8 ;
      RECT 16.8 404.4 19.8 405.6 ;
      RECT 16.8 396.3 18 405.6 ;
      RECT 14.1 396.3 24.6 397.5 ;
      RECT 7.5 -13.2 8.7 432 ;
      RECT 7.5 396.3 10.8 397.5 ;
      RECT 7.5 381.9 18 383.1 ;
      RECT 7.5 342.3 10.8 343.5 ;
      RECT 7.5 327.9 18 329.1 ;
      RECT 7.5 288.3 10.8 289.5 ;
      RECT 7.5 273.9 18 275.1 ;
      RECT 7.5 234.3 10.8 235.5 ;
      RECT 7.5 219.9 18 221.1 ;
      RECT 7.5 180.3 10.8 181.5 ;
      RECT 7.5 165.9 18 167.1 ;
      RECT 7.5 126.3 10.8 127.5 ;
      RECT 7.5 111.9 18 113.1 ;
      RECT 7.5 72.3 10.8 73.5 ;
      RECT 7.5 57.9 18 59.1 ;
      RECT 7.5 18.3 10.8 19.5 ;
      RECT 7.5 3.9 18 5.1 ;
      RECT 5.4 2.4 6.6 14.7 ;
      RECT 5.1 2.4 6.6 3.9 ;
      RECT 5.4 56.4 6.6 68.7 ;
      RECT 5.1 56.4 6.6 57.9 ;
      RECT 5.4 110.4 6.6 122.7 ;
      RECT 5.1 110.4 6.6 111.9 ;
      RECT 5.4 164.4 6.6 176.7 ;
      RECT 5.1 164.4 6.6 165.9 ;
      RECT 5.4 218.4 6.6 230.7 ;
      RECT 5.1 218.4 6.6 219.9 ;
      RECT 5.4 272.4 6.6 284.7 ;
      RECT 5.1 272.4 6.6 273.9 ;
      RECT 5.4 326.4 6.6 338.7 ;
      RECT 5.1 326.4 6.6 327.9 ;
      RECT 5.4 380.4 6.6 392.7 ;
      RECT 5.1 380.4 6.6 381.9 ;
      RECT 96 37.2 115.2 38.4 ;
      RECT 109.8 39.3 115.2 40.5 ;
      RECT 96 91.2 115.2 92.4 ;
      RECT 109.8 93.3 115.2 94.5 ;
      RECT 96 145.2 115.2 146.4 ;
      RECT 109.8 147.3 115.2 148.5 ;
      RECT 96 199.2 115.2 200.4 ;
      RECT 109.8 201.3 115.2 202.5 ;
      RECT 96 253.2 115.2 254.4 ;
      RECT 109.8 255.3 115.2 256.5 ;
      RECT 96 307.2 115.2 308.4 ;
      RECT 109.8 309.3 115.2 310.5 ;
      RECT 96 361.2 115.2 362.4 ;
      RECT 109.8 363.3 115.2 364.5 ;
      RECT 96 415.2 115.2 416.4 ;
      RECT 109.8 417.3 115.2 418.5 ;
      RECT 102.6 41.4 113.1 42.6 ;
      RECT 102.6 95.4 113.1 96.6 ;
      RECT 102.6 149.4 113.1 150.6 ;
      RECT 102.6 203.4 113.1 204.6 ;
      RECT 102.6 257.4 113.1 258.6 ;
      RECT 102.6 311.4 113.1 312.6 ;
      RECT 102.6 365.4 113.1 366.6 ;
      RECT 102.6 419.4 113.1 420.6 ;
      RECT 89.1 13.5 97.2 14.7 ;
      RECT 89.1 67.5 97.2 68.7 ;
      RECT 89.1 121.5 97.2 122.7 ;
      RECT 89.1 175.5 97.2 176.7 ;
      RECT 89.1 229.5 97.2 230.7 ;
      RECT 89.1 283.5 97.2 284.7 ;
      RECT 89.1 337.5 97.2 338.7 ;
      RECT 89.1 391.5 97.2 392.7 ;
      RECT 84.9 15.6 86.1 68.7 ;
      RECT 84.9 69.6 86.1 122.7 ;
      RECT 84.9 123.6 86.1 176.7 ;
      RECT 84.9 177.6 86.1 230.7 ;
      RECT 84.9 231.6 86.1 284.7 ;
      RECT 84.9 285.6 86.1 338.7 ;
      RECT 84.9 339.6 86.1 392.7 ;
      RECT 84.9 393.6 86.1 432 ;
      RECT 82.8 0 84 432 ;
      RECT 80.7 -5.1 81.9 432 ;
      RECT 78.6 -2.4 79.8 432 ;
      RECT 76.5 -7.8 77.7 432 ;
      RECT 74.4 -10.5 75.6 432 ;
      RECT 9.6 15.6 22.5 16.8 ;
      RECT 9.6 69.6 22.5 70.8 ;
      RECT 9.6 123.6 22.5 124.8 ;
      RECT 9.6 177.6 22.5 178.8 ;
      RECT 9.6 231.6 22.5 232.8 ;
      RECT 9.6 285.6 22.5 286.8 ;
      RECT 9.6 339.6 22.5 340.8 ;
      RECT 9.6 393.6 22.5 394.8 ;
      RECT 9.6 13.5 17.7 14.7 ;
      RECT 9.6 67.5 17.7 68.7 ;
      RECT 9.6 121.5 17.7 122.7 ;
      RECT 9.6 175.5 17.7 176.7 ;
      RECT 9.6 229.5 17.7 230.7 ;
      RECT 9.6 283.5 17.7 284.7 ;
      RECT 9.6 337.5 17.7 338.7 ;
      RECT 9.6 391.5 17.7 392.7 ;
      RECT 3 -5.1 4.2 432 ;
      RECT 0.9 -2.4 2.1 432 ;
    LAYER metal1 ;
      RECT 105 17.4 106.2 47.4 ;
      RECT 100.2 24.3 101.4 33.6 ;
      RECT 87.3 24.3 153 29.7 ;
      RECT 139.2 20.4 140.7 29.7 ;
      RECT 131.4 20.4 132.6 29.7 ;
      RECT 126.3 20.4 127.8 29.7 ;
      RECT 118.5 20.4 119.7 29.7 ;
      RECT 112.2 20.4 113.4 29.7 ;
      RECT 91.2 20.4 92.4 29.7 ;
      RECT 139.2 51.3 140.7 63.6 ;
      RECT 131.4 51.3 132.6 63.6 ;
      RECT 126.3 51.3 127.8 63.6 ;
      RECT 118.5 51.3 119.7 63.6 ;
      RECT 112.2 51.3 113.4 63.6 ;
      RECT 109.8 51.3 111 63.6 ;
      RECT 105 51.3 106.2 63.6 ;
      RECT 91.2 51.3 92.4 63.6 ;
      RECT 59.7 51.3 61.2 63.6 ;
      RECT 51.9 51.3 53.1 63.6 ;
      RECT 46.8 51.3 48.3 63.6 ;
      RECT 39 44.4 40.2 63.6 ;
      RECT 32.7 44.4 33.9 63.6 ;
      RECT 30.3 51.3 31.5 63.6 ;
      RECT 28.8 51.3 153 56.7 ;
      RECT 100.2 44.4 101.4 56.7 ;
      RECT 66 44.4 67.2 56.7 ;
      RECT 61.2 44.4 62.4 56.7 ;
      RECT 53.4 44.4 54.6 56.7 ;
      RECT 43.8 44.4 45 56.7 ;
      RECT 105 71.4 106.2 101.4 ;
      RECT 16.5 78.3 17.7 101.4 ;
      RECT 100.2 78.3 101.4 87.6 ;
      RECT 66 78.3 67.2 87.6 ;
      RECT 61.2 78.3 62.4 87.6 ;
      RECT 53.4 78.3 54.6 87.6 ;
      RECT 43.8 78.3 45 87.6 ;
      RECT 39 74.4 40.2 87.6 ;
      RECT 32.7 74.4 33.9 87.6 ;
      RECT 25.5 71.4 26.7 87.6 ;
      RECT 20.7 78.3 21.9 87.6 ;
      RECT 0 78.3 153 83.7 ;
      RECT 139.2 74.4 140.7 83.7 ;
      RECT 131.4 74.4 132.6 83.7 ;
      RECT 126.3 74.4 127.8 83.7 ;
      RECT 118.5 74.4 119.7 83.7 ;
      RECT 112.2 74.4 113.4 83.7 ;
      RECT 91.2 74.4 92.4 83.7 ;
      RECT 59.7 74.4 61.2 83.7 ;
      RECT 51.9 74.4 53.1 83.7 ;
      RECT 46.8 74.4 48.3 83.7 ;
      RECT 11.7 74.4 12.9 83.7 ;
      RECT 7.5 69.6 8.7 83.7 ;
      RECT 6.9 69.6 10.8 70.8 ;
      RECT 139.2 105.3 140.7 117.6 ;
      RECT 131.4 105.3 132.6 117.6 ;
      RECT 126.3 105.3 127.8 117.6 ;
      RECT 118.5 105.3 119.7 117.6 ;
      RECT 112.2 105.3 113.4 117.6 ;
      RECT 109.8 105.3 111 117.6 ;
      RECT 105 105.3 106.2 117.6 ;
      RECT 91.2 105.3 92.4 117.6 ;
      RECT 59.7 105.3 61.2 117.6 ;
      RECT 51.9 105.3 53.1 117.6 ;
      RECT 46.8 105.3 48.3 117.6 ;
      RECT 39 98.4 40.2 117.6 ;
      RECT 32.7 98.4 33.9 117.6 ;
      RECT 30.3 105.3 31.5 117.6 ;
      RECT 28.8 105.3 153 110.7 ;
      RECT 100.2 98.4 101.4 110.7 ;
      RECT 66 98.4 67.2 110.7 ;
      RECT 61.2 98.4 62.4 110.7 ;
      RECT 53.4 98.4 54.6 110.7 ;
      RECT 43.8 98.4 45 110.7 ;
      RECT 105 125.4 106.2 155.4 ;
      RECT 16.5 132.3 17.7 155.4 ;
      RECT 100.2 132.3 101.4 141.6 ;
      RECT 66 132.3 67.2 141.6 ;
      RECT 61.2 132.3 62.4 141.6 ;
      RECT 53.4 132.3 54.6 141.6 ;
      RECT 43.8 132.3 45 141.6 ;
      RECT 39 128.4 40.2 141.6 ;
      RECT 32.7 128.4 33.9 141.6 ;
      RECT 25.5 125.4 26.7 141.6 ;
      RECT 20.7 132.3 21.9 141.6 ;
      RECT 0 132.3 153 137.7 ;
      RECT 139.2 128.4 140.7 137.7 ;
      RECT 131.4 128.4 132.6 137.7 ;
      RECT 126.3 128.4 127.8 137.7 ;
      RECT 118.5 128.4 119.7 137.7 ;
      RECT 112.2 128.4 113.4 137.7 ;
      RECT 91.2 128.4 92.4 137.7 ;
      RECT 59.7 128.4 61.2 137.7 ;
      RECT 51.9 128.4 53.1 137.7 ;
      RECT 46.8 128.4 48.3 137.7 ;
      RECT 11.7 128.4 12.9 137.7 ;
      RECT 7.5 123.6 8.7 137.7 ;
      RECT 6.9 123.6 10.8 124.8 ;
      RECT 139.2 159.3 140.7 171.6 ;
      RECT 131.4 159.3 132.6 171.6 ;
      RECT 126.3 159.3 127.8 171.6 ;
      RECT 118.5 159.3 119.7 171.6 ;
      RECT 112.2 159.3 113.4 171.6 ;
      RECT 109.8 159.3 111 171.6 ;
      RECT 105 159.3 106.2 171.6 ;
      RECT 91.2 159.3 92.4 171.6 ;
      RECT 59.7 159.3 61.2 171.6 ;
      RECT 51.9 159.3 53.1 171.6 ;
      RECT 46.8 159.3 48.3 171.6 ;
      RECT 39 152.4 40.2 171.6 ;
      RECT 32.7 152.4 33.9 171.6 ;
      RECT 30.3 159.3 31.5 171.6 ;
      RECT 28.8 159.3 153 164.7 ;
      RECT 100.2 152.4 101.4 164.7 ;
      RECT 66 152.4 67.2 164.7 ;
      RECT 61.2 152.4 62.4 164.7 ;
      RECT 53.4 152.4 54.6 164.7 ;
      RECT 43.8 152.4 45 164.7 ;
      RECT 105 179.4 106.2 209.4 ;
      RECT 16.5 186.3 17.7 209.4 ;
      RECT 100.2 186.3 101.4 195.6 ;
      RECT 66 186.3 67.2 195.6 ;
      RECT 61.2 186.3 62.4 195.6 ;
      RECT 53.4 186.3 54.6 195.6 ;
      RECT 43.8 186.3 45 195.6 ;
      RECT 39 182.4 40.2 195.6 ;
      RECT 32.7 182.4 33.9 195.6 ;
      RECT 25.5 179.4 26.7 195.6 ;
      RECT 20.7 186.3 21.9 195.6 ;
      RECT 0 186.3 153 191.7 ;
      RECT 139.2 182.4 140.7 191.7 ;
      RECT 131.4 182.4 132.6 191.7 ;
      RECT 126.3 182.4 127.8 191.7 ;
      RECT 118.5 182.4 119.7 191.7 ;
      RECT 112.2 182.4 113.4 191.7 ;
      RECT 91.2 182.4 92.4 191.7 ;
      RECT 59.7 182.4 61.2 191.7 ;
      RECT 51.9 182.4 53.1 191.7 ;
      RECT 46.8 182.4 48.3 191.7 ;
      RECT 11.7 182.4 12.9 191.7 ;
      RECT 7.5 177.6 8.7 191.7 ;
      RECT 6.9 177.6 10.8 178.8 ;
      RECT 139.2 213.3 140.7 225.6 ;
      RECT 131.4 213.3 132.6 225.6 ;
      RECT 126.3 213.3 127.8 225.6 ;
      RECT 118.5 213.3 119.7 225.6 ;
      RECT 112.2 213.3 113.4 225.6 ;
      RECT 109.8 213.3 111 225.6 ;
      RECT 105 213.3 106.2 225.6 ;
      RECT 91.2 213.3 92.4 225.6 ;
      RECT 59.7 213.3 61.2 225.6 ;
      RECT 51.9 213.3 53.1 225.6 ;
      RECT 46.8 213.3 48.3 225.6 ;
      RECT 39 206.4 40.2 225.6 ;
      RECT 32.7 206.4 33.9 225.6 ;
      RECT 30.3 213.3 31.5 225.6 ;
      RECT 28.8 213.3 153 218.7 ;
      RECT 100.2 206.4 101.4 218.7 ;
      RECT 66 206.4 67.2 218.7 ;
      RECT 61.2 206.4 62.4 218.7 ;
      RECT 53.4 206.4 54.6 218.7 ;
      RECT 43.8 206.4 45 218.7 ;
      RECT 105 233.4 106.2 263.4 ;
      RECT 16.5 240.3 17.7 263.4 ;
      RECT 100.2 240.3 101.4 249.6 ;
      RECT 66 240.3 67.2 249.6 ;
      RECT 61.2 240.3 62.4 249.6 ;
      RECT 53.4 240.3 54.6 249.6 ;
      RECT 43.8 240.3 45 249.6 ;
      RECT 39 236.4 40.2 249.6 ;
      RECT 32.7 236.4 33.9 249.6 ;
      RECT 25.5 233.4 26.7 249.6 ;
      RECT 20.7 240.3 21.9 249.6 ;
      RECT 0 240.3 153 245.7 ;
      RECT 139.2 236.4 140.7 245.7 ;
      RECT 131.4 236.4 132.6 245.7 ;
      RECT 126.3 236.4 127.8 245.7 ;
      RECT 118.5 236.4 119.7 245.7 ;
      RECT 112.2 236.4 113.4 245.7 ;
      RECT 91.2 236.4 92.4 245.7 ;
      RECT 59.7 236.4 61.2 245.7 ;
      RECT 51.9 236.4 53.1 245.7 ;
      RECT 46.8 236.4 48.3 245.7 ;
      RECT 11.7 236.4 12.9 245.7 ;
      RECT 7.5 231.6 8.7 245.7 ;
      RECT 6.9 231.6 10.8 232.8 ;
      RECT 139.2 267.3 140.7 279.6 ;
      RECT 131.4 267.3 132.6 279.6 ;
      RECT 126.3 267.3 127.8 279.6 ;
      RECT 118.5 267.3 119.7 279.6 ;
      RECT 112.2 267.3 113.4 279.6 ;
      RECT 109.8 267.3 111 279.6 ;
      RECT 105 267.3 106.2 279.6 ;
      RECT 91.2 267.3 92.4 279.6 ;
      RECT 59.7 267.3 61.2 279.6 ;
      RECT 51.9 267.3 53.1 279.6 ;
      RECT 46.8 267.3 48.3 279.6 ;
      RECT 39 260.4 40.2 279.6 ;
      RECT 32.7 260.4 33.9 279.6 ;
      RECT 30.3 267.3 31.5 279.6 ;
      RECT 28.8 267.3 153 272.7 ;
      RECT 100.2 260.4 101.4 272.7 ;
      RECT 66 260.4 67.2 272.7 ;
      RECT 61.2 260.4 62.4 272.7 ;
      RECT 53.4 260.4 54.6 272.7 ;
      RECT 43.8 260.4 45 272.7 ;
      RECT 105 287.4 106.2 317.4 ;
      RECT 16.5 294.3 17.7 317.4 ;
      RECT 100.2 294.3 101.4 303.6 ;
      RECT 66 294.3 67.2 303.6 ;
      RECT 61.2 294.3 62.4 303.6 ;
      RECT 53.4 294.3 54.6 303.6 ;
      RECT 43.8 294.3 45 303.6 ;
      RECT 39 290.4 40.2 303.6 ;
      RECT 32.7 290.4 33.9 303.6 ;
      RECT 25.5 287.4 26.7 303.6 ;
      RECT 20.7 294.3 21.9 303.6 ;
      RECT 0 294.3 153 299.7 ;
      RECT 139.2 290.4 140.7 299.7 ;
      RECT 131.4 290.4 132.6 299.7 ;
      RECT 126.3 290.4 127.8 299.7 ;
      RECT 118.5 290.4 119.7 299.7 ;
      RECT 112.2 290.4 113.4 299.7 ;
      RECT 91.2 290.4 92.4 299.7 ;
      RECT 59.7 290.4 61.2 299.7 ;
      RECT 51.9 290.4 53.1 299.7 ;
      RECT 46.8 290.4 48.3 299.7 ;
      RECT 11.7 290.4 12.9 299.7 ;
      RECT 7.5 285.6 8.7 299.7 ;
      RECT 6.9 285.6 10.8 286.8 ;
      RECT 139.2 321.3 140.7 333.6 ;
      RECT 131.4 321.3 132.6 333.6 ;
      RECT 126.3 321.3 127.8 333.6 ;
      RECT 118.5 321.3 119.7 333.6 ;
      RECT 112.2 321.3 113.4 333.6 ;
      RECT 109.8 321.3 111 333.6 ;
      RECT 105 321.3 106.2 333.6 ;
      RECT 91.2 321.3 92.4 333.6 ;
      RECT 59.7 321.3 61.2 333.6 ;
      RECT 51.9 321.3 53.1 333.6 ;
      RECT 46.8 321.3 48.3 333.6 ;
      RECT 39 314.4 40.2 333.6 ;
      RECT 32.7 314.4 33.9 333.6 ;
      RECT 30.3 321.3 31.5 333.6 ;
      RECT 28.8 321.3 153 326.7 ;
      RECT 100.2 314.4 101.4 326.7 ;
      RECT 66 314.4 67.2 326.7 ;
      RECT 61.2 314.4 62.4 326.7 ;
      RECT 53.4 314.4 54.6 326.7 ;
      RECT 43.8 314.4 45 326.7 ;
      RECT 105 341.4 106.2 371.4 ;
      RECT 16.5 348.3 17.7 371.4 ;
      RECT 100.2 348.3 101.4 357.6 ;
      RECT 66 348.3 67.2 357.6 ;
      RECT 61.2 348.3 62.4 357.6 ;
      RECT 53.4 348.3 54.6 357.6 ;
      RECT 43.8 348.3 45 357.6 ;
      RECT 39 344.4 40.2 357.6 ;
      RECT 32.7 344.4 33.9 357.6 ;
      RECT 25.5 341.4 26.7 357.6 ;
      RECT 20.7 348.3 21.9 357.6 ;
      RECT 0 348.3 153 353.7 ;
      RECT 139.2 344.4 140.7 353.7 ;
      RECT 131.4 344.4 132.6 353.7 ;
      RECT 126.3 344.4 127.8 353.7 ;
      RECT 118.5 344.4 119.7 353.7 ;
      RECT 112.2 344.4 113.4 353.7 ;
      RECT 91.2 344.4 92.4 353.7 ;
      RECT 59.7 344.4 61.2 353.7 ;
      RECT 51.9 344.4 53.1 353.7 ;
      RECT 46.8 344.4 48.3 353.7 ;
      RECT 11.7 344.4 12.9 353.7 ;
      RECT 7.5 339.6 8.7 353.7 ;
      RECT 6.9 339.6 10.8 340.8 ;
      RECT 139.2 375.3 140.7 387.6 ;
      RECT 131.4 375.3 132.6 387.6 ;
      RECT 126.3 375.3 127.8 387.6 ;
      RECT 118.5 375.3 119.7 387.6 ;
      RECT 112.2 375.3 113.4 387.6 ;
      RECT 109.8 375.3 111 387.6 ;
      RECT 105 375.3 106.2 387.6 ;
      RECT 91.2 375.3 92.4 387.6 ;
      RECT 59.7 375.3 61.2 387.6 ;
      RECT 51.9 375.3 53.1 387.6 ;
      RECT 46.8 375.3 48.3 387.6 ;
      RECT 39 368.4 40.2 387.6 ;
      RECT 32.7 368.4 33.9 387.6 ;
      RECT 30.3 375.3 31.5 387.6 ;
      RECT 28.8 375.3 153 380.7 ;
      RECT 100.2 368.4 101.4 380.7 ;
      RECT 66 368.4 67.2 380.7 ;
      RECT 61.2 368.4 62.4 380.7 ;
      RECT 53.4 368.4 54.6 380.7 ;
      RECT 43.8 368.4 45 380.7 ;
      RECT 105 395.4 106.2 425.4 ;
      RECT 100.2 402.3 101.4 411.6 ;
      RECT 87.3 402.3 153 407.7 ;
      RECT 139.2 398.4 140.7 407.7 ;
      RECT 131.4 398.4 132.6 407.7 ;
      RECT 126.3 398.4 127.8 407.7 ;
      RECT 118.5 398.4 119.7 407.7 ;
      RECT 112.2 398.4 113.4 407.7 ;
      RECT 91.2 398.4 92.4 407.7 ;
      RECT 143.4 15.9 144.6 23.4 ;
      RECT 138.6 18.3 144.6 19.5 ;
      RECT 143.4 3.6 143.7 23.4 ;
      RECT 143.4 3.6 144.6 12.6 ;
      RECT 143.4 69.9 144.6 77.4 ;
      RECT 138.6 72.3 144.6 73.5 ;
      RECT 143.4 57.6 143.7 77.4 ;
      RECT 143.4 57.6 144.6 66.6 ;
      RECT 143.4 123.9 144.6 131.4 ;
      RECT 138.6 126.3 144.6 127.5 ;
      RECT 143.4 111.6 143.7 131.4 ;
      RECT 143.4 111.6 144.6 120.6 ;
      RECT 143.4 177.9 144.6 185.4 ;
      RECT 138.6 180.3 144.6 181.5 ;
      RECT 143.4 165.6 143.7 185.4 ;
      RECT 143.4 165.6 144.6 174.6 ;
      RECT 143.4 231.9 144.6 239.4 ;
      RECT 138.6 234.3 144.6 235.5 ;
      RECT 143.4 219.6 143.7 239.4 ;
      RECT 143.4 219.6 144.6 228.6 ;
      RECT 143.4 285.9 144.6 293.4 ;
      RECT 138.6 288.3 144.6 289.5 ;
      RECT 143.4 273.6 143.7 293.4 ;
      RECT 143.4 273.6 144.6 282.6 ;
      RECT 143.4 339.9 144.6 347.4 ;
      RECT 138.6 342.3 144.6 343.5 ;
      RECT 143.4 327.6 143.7 347.4 ;
      RECT 143.4 327.6 144.6 336.6 ;
      RECT 143.4 393.9 144.6 401.4 ;
      RECT 138.6 396.3 144.6 397.5 ;
      RECT 143.4 381.6 143.7 401.4 ;
      RECT 143.4 381.6 144.6 390.6 ;
      RECT 135.3 20.4 136.5 23.4 ;
      RECT 135.6 16.5 136.5 23.4 ;
      RECT 135.6 16.5 141.3 17.4 ;
      RECT 140.1 10.5 141.3 17.4 ;
      RECT 135.6 10.5 141.3 11.7 ;
      RECT 135.6 3.6 136.5 11.7 ;
      RECT 135.3 3.6 136.5 9.6 ;
      RECT 135.3 74.4 136.5 77.4 ;
      RECT 135.6 70.5 136.5 77.4 ;
      RECT 135.6 70.5 141.3 71.4 ;
      RECT 140.1 64.5 141.3 71.4 ;
      RECT 135.6 64.5 141.3 65.7 ;
      RECT 135.6 57.6 136.5 65.7 ;
      RECT 135.3 57.6 136.5 63.6 ;
      RECT 135.3 128.4 136.5 131.4 ;
      RECT 135.6 124.5 136.5 131.4 ;
      RECT 135.6 124.5 141.3 125.4 ;
      RECT 140.1 118.5 141.3 125.4 ;
      RECT 135.6 118.5 141.3 119.7 ;
      RECT 135.6 111.6 136.5 119.7 ;
      RECT 135.3 111.6 136.5 117.6 ;
      RECT 135.3 182.4 136.5 185.4 ;
      RECT 135.6 178.5 136.5 185.4 ;
      RECT 135.6 178.5 141.3 179.4 ;
      RECT 140.1 172.5 141.3 179.4 ;
      RECT 135.6 172.5 141.3 173.7 ;
      RECT 135.6 165.6 136.5 173.7 ;
      RECT 135.3 165.6 136.5 171.6 ;
      RECT 135.3 236.4 136.5 239.4 ;
      RECT 135.6 232.5 136.5 239.4 ;
      RECT 135.6 232.5 141.3 233.4 ;
      RECT 140.1 226.5 141.3 233.4 ;
      RECT 135.6 226.5 141.3 227.7 ;
      RECT 135.6 219.6 136.5 227.7 ;
      RECT 135.3 219.6 136.5 225.6 ;
      RECT 135.3 290.4 136.5 293.4 ;
      RECT 135.6 286.5 136.5 293.4 ;
      RECT 135.6 286.5 141.3 287.4 ;
      RECT 140.1 280.5 141.3 287.4 ;
      RECT 135.6 280.5 141.3 281.7 ;
      RECT 135.6 273.6 136.5 281.7 ;
      RECT 135.3 273.6 136.5 279.6 ;
      RECT 135.3 344.4 136.5 347.4 ;
      RECT 135.6 340.5 136.5 347.4 ;
      RECT 135.6 340.5 141.3 341.4 ;
      RECT 140.1 334.5 141.3 341.4 ;
      RECT 135.6 334.5 141.3 335.7 ;
      RECT 135.6 327.6 136.5 335.7 ;
      RECT 135.3 327.6 136.5 333.6 ;
      RECT 135.3 398.4 136.5 401.4 ;
      RECT 135.6 394.5 136.5 401.4 ;
      RECT 135.6 394.5 141.3 395.4 ;
      RECT 140.1 388.5 141.3 395.4 ;
      RECT 135.6 388.5 141.3 389.7 ;
      RECT 135.6 381.6 136.5 389.7 ;
      RECT 135.3 381.6 136.5 387.6 ;
      RECT 129 18.3 130.2 23.4 ;
      RECT 129.3 3.6 130.2 23.4 ;
      RECT 125.7 18.3 130.2 19.5 ;
      RECT 129.3 13.5 131.1 14.7 ;
      RECT 129 3.6 130.2 9.6 ;
      RECT 129 72.3 130.2 77.4 ;
      RECT 129.3 57.6 130.2 77.4 ;
      RECT 125.7 72.3 130.2 73.5 ;
      RECT 129.3 67.5 131.1 68.7 ;
      RECT 129 57.6 130.2 63.6 ;
      RECT 129 126.3 130.2 131.4 ;
      RECT 129.3 111.6 130.2 131.4 ;
      RECT 125.7 126.3 130.2 127.5 ;
      RECT 129.3 121.5 131.1 122.7 ;
      RECT 129 111.6 130.2 117.6 ;
      RECT 129 180.3 130.2 185.4 ;
      RECT 129.3 165.6 130.2 185.4 ;
      RECT 125.7 180.3 130.2 181.5 ;
      RECT 129.3 175.5 131.1 176.7 ;
      RECT 129 165.6 130.2 171.6 ;
      RECT 129 234.3 130.2 239.4 ;
      RECT 129.3 219.6 130.2 239.4 ;
      RECT 125.7 234.3 130.2 235.5 ;
      RECT 129.3 229.5 131.1 230.7 ;
      RECT 129 219.6 130.2 225.6 ;
      RECT 129 288.3 130.2 293.4 ;
      RECT 129.3 273.6 130.2 293.4 ;
      RECT 125.7 288.3 130.2 289.5 ;
      RECT 129.3 283.5 131.1 284.7 ;
      RECT 129 273.6 130.2 279.6 ;
      RECT 129 342.3 130.2 347.4 ;
      RECT 129.3 327.6 130.2 347.4 ;
      RECT 125.7 342.3 130.2 343.5 ;
      RECT 129.3 337.5 131.1 338.7 ;
      RECT 129 327.6 130.2 333.6 ;
      RECT 129 396.3 130.2 401.4 ;
      RECT 129.3 381.6 130.2 401.4 ;
      RECT 125.7 396.3 130.2 397.5 ;
      RECT 129.3 391.5 131.1 392.7 ;
      RECT 129 381.6 130.2 387.6 ;
      RECT 122.4 20.4 123.6 23.4 ;
      RECT 122.7 16.5 123.6 23.4 ;
      RECT 122.7 16.5 128.4 17.4 ;
      RECT 127.2 10.5 128.4 17.4 ;
      RECT 122.7 10.5 128.4 11.7 ;
      RECT 122.7 3.6 123.6 11.7 ;
      RECT 122.4 3.6 123.6 9.6 ;
      RECT 122.4 74.4 123.6 77.4 ;
      RECT 122.7 70.5 123.6 77.4 ;
      RECT 122.7 70.5 128.4 71.4 ;
      RECT 127.2 64.5 128.4 71.4 ;
      RECT 122.7 64.5 128.4 65.7 ;
      RECT 122.7 57.6 123.6 65.7 ;
      RECT 122.4 57.6 123.6 63.6 ;
      RECT 122.4 128.4 123.6 131.4 ;
      RECT 122.7 124.5 123.6 131.4 ;
      RECT 122.7 124.5 128.4 125.4 ;
      RECT 127.2 118.5 128.4 125.4 ;
      RECT 122.7 118.5 128.4 119.7 ;
      RECT 122.7 111.6 123.6 119.7 ;
      RECT 122.4 111.6 123.6 117.6 ;
      RECT 122.4 182.4 123.6 185.4 ;
      RECT 122.7 178.5 123.6 185.4 ;
      RECT 122.7 178.5 128.4 179.4 ;
      RECT 127.2 172.5 128.4 179.4 ;
      RECT 122.7 172.5 128.4 173.7 ;
      RECT 122.7 165.6 123.6 173.7 ;
      RECT 122.4 165.6 123.6 171.6 ;
      RECT 122.4 236.4 123.6 239.4 ;
      RECT 122.7 232.5 123.6 239.4 ;
      RECT 122.7 232.5 128.4 233.4 ;
      RECT 127.2 226.5 128.4 233.4 ;
      RECT 122.7 226.5 128.4 227.7 ;
      RECT 122.7 219.6 123.6 227.7 ;
      RECT 122.4 219.6 123.6 225.6 ;
      RECT 122.4 290.4 123.6 293.4 ;
      RECT 122.7 286.5 123.6 293.4 ;
      RECT 122.7 286.5 128.4 287.4 ;
      RECT 127.2 280.5 128.4 287.4 ;
      RECT 122.7 280.5 128.4 281.7 ;
      RECT 122.7 273.6 123.6 281.7 ;
      RECT 122.4 273.6 123.6 279.6 ;
      RECT 122.4 344.4 123.6 347.4 ;
      RECT 122.7 340.5 123.6 347.4 ;
      RECT 122.7 340.5 128.4 341.4 ;
      RECT 127.2 334.5 128.4 341.4 ;
      RECT 122.7 334.5 128.4 335.7 ;
      RECT 122.7 327.6 123.6 335.7 ;
      RECT 122.4 327.6 123.6 333.6 ;
      RECT 122.4 398.4 123.6 401.4 ;
      RECT 122.7 394.5 123.6 401.4 ;
      RECT 122.7 394.5 128.4 395.4 ;
      RECT 127.2 388.5 128.4 395.4 ;
      RECT 122.7 388.5 128.4 389.7 ;
      RECT 122.7 381.6 123.6 389.7 ;
      RECT 122.4 381.6 123.6 387.6 ;
      RECT 116.1 3.6 117.3 23.4 ;
      RECT 120.6 10.5 121.8 12.9 ;
      RECT 116.1 10.5 121.8 11.7 ;
      RECT 116.1 57.6 117.3 77.4 ;
      RECT 120.6 64.5 121.8 66.9 ;
      RECT 116.1 64.5 121.8 65.7 ;
      RECT 116.1 111.6 117.3 131.4 ;
      RECT 120.6 118.5 121.8 120.9 ;
      RECT 116.1 118.5 121.8 119.7 ;
      RECT 116.1 165.6 117.3 185.4 ;
      RECT 120.6 172.5 121.8 174.9 ;
      RECT 116.1 172.5 121.8 173.7 ;
      RECT 116.1 219.6 117.3 239.4 ;
      RECT 120.6 226.5 121.8 228.9 ;
      RECT 116.1 226.5 121.8 227.7 ;
      RECT 116.1 273.6 117.3 293.4 ;
      RECT 120.6 280.5 121.8 282.9 ;
      RECT 116.1 280.5 121.8 281.7 ;
      RECT 116.1 327.6 117.3 347.4 ;
      RECT 120.6 334.5 121.8 336.9 ;
      RECT 116.1 334.5 121.8 335.7 ;
      RECT 116.1 381.6 117.3 401.4 ;
      RECT 120.6 388.5 121.8 390.9 ;
      RECT 116.1 388.5 121.8 389.7 ;
      RECT 108.9 17.4 110.1 23.4 ;
      RECT 113.7 17.1 114.9 19.5 ;
      RECT 108.9 17.4 114.9 18.3 ;
      RECT 110.4 17.1 114.9 18.3 ;
      RECT 110.4 10.5 111.3 18.3 ;
      RECT 107.7 10.5 111.3 11.4 ;
      RECT 107.7 3.6 108.6 11.4 ;
      RECT 107.4 3.6 108.6 9.6 ;
      RECT 108.9 71.4 110.1 77.4 ;
      RECT 113.7 71.1 114.9 73.5 ;
      RECT 108.9 71.4 114.9 72.3 ;
      RECT 110.4 71.1 114.9 72.3 ;
      RECT 110.4 64.5 111.3 72.3 ;
      RECT 107.7 64.5 111.3 65.4 ;
      RECT 107.7 57.6 108.6 65.4 ;
      RECT 107.4 57.6 108.6 63.6 ;
      RECT 108.9 125.4 110.1 131.4 ;
      RECT 113.7 125.1 114.9 127.5 ;
      RECT 108.9 125.4 114.9 126.3 ;
      RECT 110.4 125.1 114.9 126.3 ;
      RECT 110.4 118.5 111.3 126.3 ;
      RECT 107.7 118.5 111.3 119.4 ;
      RECT 107.7 111.6 108.6 119.4 ;
      RECT 107.4 111.6 108.6 117.6 ;
      RECT 108.9 179.4 110.1 185.4 ;
      RECT 113.7 179.1 114.9 181.5 ;
      RECT 108.9 179.4 114.9 180.3 ;
      RECT 110.4 179.1 114.9 180.3 ;
      RECT 110.4 172.5 111.3 180.3 ;
      RECT 107.7 172.5 111.3 173.4 ;
      RECT 107.7 165.6 108.6 173.4 ;
      RECT 107.4 165.6 108.6 171.6 ;
      RECT 108.9 233.4 110.1 239.4 ;
      RECT 113.7 233.1 114.9 235.5 ;
      RECT 108.9 233.4 114.9 234.3 ;
      RECT 110.4 233.1 114.9 234.3 ;
      RECT 110.4 226.5 111.3 234.3 ;
      RECT 107.7 226.5 111.3 227.4 ;
      RECT 107.7 219.6 108.6 227.4 ;
      RECT 107.4 219.6 108.6 225.6 ;
      RECT 108.9 287.4 110.1 293.4 ;
      RECT 113.7 287.1 114.9 289.5 ;
      RECT 108.9 287.4 114.9 288.3 ;
      RECT 110.4 287.1 114.9 288.3 ;
      RECT 110.4 280.5 111.3 288.3 ;
      RECT 107.7 280.5 111.3 281.4 ;
      RECT 107.7 273.6 108.6 281.4 ;
      RECT 107.4 273.6 108.6 279.6 ;
      RECT 108.9 341.4 110.1 347.4 ;
      RECT 113.7 341.1 114.9 343.5 ;
      RECT 108.9 341.4 114.9 342.3 ;
      RECT 110.4 341.1 114.9 342.3 ;
      RECT 110.4 334.5 111.3 342.3 ;
      RECT 107.7 334.5 111.3 335.4 ;
      RECT 107.7 327.6 108.6 335.4 ;
      RECT 107.4 327.6 108.6 333.6 ;
      RECT 108.9 395.4 110.1 401.4 ;
      RECT 113.7 395.1 114.9 397.5 ;
      RECT 108.9 395.4 114.9 396.3 ;
      RECT 110.4 395.1 114.9 396.3 ;
      RECT 110.4 388.5 111.3 396.3 ;
      RECT 107.7 388.5 111.3 389.4 ;
      RECT 107.7 381.6 108.6 389.4 ;
      RECT 107.4 381.6 108.6 387.6 ;
      RECT 91.2 30.6 92.4 47.4 ;
      RECT 86.4 30.6 92.4 31.8 ;
      RECT 91.2 84.6 92.4 101.4 ;
      RECT 86.4 84.6 92.4 85.8 ;
      RECT 91.2 138.6 92.4 155.4 ;
      RECT 86.4 138.6 92.4 139.8 ;
      RECT 91.2 192.6 92.4 209.4 ;
      RECT 86.4 192.6 92.4 193.8 ;
      RECT 91.2 246.6 92.4 263.4 ;
      RECT 86.4 246.6 92.4 247.8 ;
      RECT 91.2 300.6 92.4 317.4 ;
      RECT 86.4 300.6 92.4 301.8 ;
      RECT 91.2 354.6 92.4 371.4 ;
      RECT 86.4 354.6 92.4 355.8 ;
      RECT 91.2 408.6 92.4 425.4 ;
      RECT 82.8 419.4 90.3 420.6 ;
      RECT 89.1 408.6 90.3 420.6 ;
      RECT 86.4 408.6 92.4 409.8 ;
      RECT 68.4 30.6 69.6 50.4 ;
      RECT 68.4 34.5 70.8 35.7 ;
      RECT 68.4 84.6 69.6 104.4 ;
      RECT 68.4 88.5 70.8 89.7 ;
      RECT 68.4 138.6 69.6 158.4 ;
      RECT 68.4 142.5 70.8 143.7 ;
      RECT 68.4 192.6 69.6 212.4 ;
      RECT 68.4 196.5 70.8 197.7 ;
      RECT 68.4 246.6 69.6 266.4 ;
      RECT 68.4 250.5 70.8 251.7 ;
      RECT 68.4 300.6 69.6 320.4 ;
      RECT 68.4 304.5 70.8 305.7 ;
      RECT 68.4 354.6 69.6 374.4 ;
      RECT 68.4 358.5 70.8 359.7 ;
      RECT 68.4 408.6 69.6 428.4 ;
      RECT 68.4 412.5 70.8 413.7 ;
      RECT 28.8 429.3 70.2 430.2 ;
      RECT 66 422.4 67.2 430.2 ;
      RECT 61.2 422.4 62.4 430.2 ;
      RECT 53.4 422.4 54.6 430.2 ;
      RECT 43.8 422.4 45 430.2 ;
      RECT 39 422.4 40.2 430.2 ;
      RECT 32.7 422.4 33.9 430.2 ;
      RECT 58.8 44.4 60 50.4 ;
      RECT 59.1 30.6 60 50.4 ;
      RECT 51 44.4 52.2 50.4 ;
      RECT 51 30.6 51.9 50.4 ;
      RECT 51 35.7 60 36.6 ;
      RECT 59.1 34.5 62.4 35.7 ;
      RECT 58.8 30.6 60 33.6 ;
      RECT 51 30.6 52.2 33.6 ;
      RECT 58.8 98.4 60 104.4 ;
      RECT 59.1 84.6 60 104.4 ;
      RECT 51 98.4 52.2 104.4 ;
      RECT 51 84.6 51.9 104.4 ;
      RECT 51 89.7 60 90.6 ;
      RECT 59.1 88.5 62.4 89.7 ;
      RECT 58.8 84.6 60 87.6 ;
      RECT 51 84.6 52.2 87.6 ;
      RECT 58.8 152.4 60 158.4 ;
      RECT 59.1 138.6 60 158.4 ;
      RECT 51 152.4 52.2 158.4 ;
      RECT 51 138.6 51.9 158.4 ;
      RECT 51 143.7 60 144.6 ;
      RECT 59.1 142.5 62.4 143.7 ;
      RECT 58.8 138.6 60 141.6 ;
      RECT 51 138.6 52.2 141.6 ;
      RECT 58.8 206.4 60 212.4 ;
      RECT 59.1 192.6 60 212.4 ;
      RECT 51 206.4 52.2 212.4 ;
      RECT 51 192.6 51.9 212.4 ;
      RECT 51 197.7 60 198.6 ;
      RECT 59.1 196.5 62.4 197.7 ;
      RECT 58.8 192.6 60 195.6 ;
      RECT 51 192.6 52.2 195.6 ;
      RECT 58.8 260.4 60 266.4 ;
      RECT 59.1 246.6 60 266.4 ;
      RECT 51 260.4 52.2 266.4 ;
      RECT 51 246.6 51.9 266.4 ;
      RECT 51 251.7 60 252.6 ;
      RECT 59.1 250.5 62.4 251.7 ;
      RECT 58.8 246.6 60 249.6 ;
      RECT 51 246.6 52.2 249.6 ;
      RECT 58.8 314.4 60 320.4 ;
      RECT 59.1 300.6 60 320.4 ;
      RECT 51 314.4 52.2 320.4 ;
      RECT 51 300.6 51.9 320.4 ;
      RECT 51 305.7 60 306.6 ;
      RECT 59.1 304.5 62.4 305.7 ;
      RECT 58.8 300.6 60 303.6 ;
      RECT 51 300.6 52.2 303.6 ;
      RECT 58.8 368.4 60 374.4 ;
      RECT 59.1 354.6 60 374.4 ;
      RECT 51 368.4 52.2 374.4 ;
      RECT 51 354.6 51.9 374.4 ;
      RECT 51 359.7 60 360.6 ;
      RECT 59.1 358.5 62.4 359.7 ;
      RECT 58.8 354.6 60 357.6 ;
      RECT 51 354.6 52.2 357.6 ;
      RECT 58.8 422.4 60 428.4 ;
      RECT 59.1 408.6 60 428.4 ;
      RECT 51 422.4 52.2 428.4 ;
      RECT 51 408.6 51.9 428.4 ;
      RECT 51 413.7 60 414.6 ;
      RECT 59.1 412.5 62.4 413.7 ;
      RECT 58.8 408.6 60 411.6 ;
      RECT 51 408.6 52.2 411.6 ;
      RECT 55.8 20.4 57 23.4 ;
      RECT 56.1 16.5 57 23.4 ;
      RECT 56.1 16.5 61.8 17.4 ;
      RECT 60.6 10.5 61.8 17.4 ;
      RECT 56.1 10.5 61.8 11.7 ;
      RECT 56.1 3.6 57 11.7 ;
      RECT 55.8 3.6 57 9.6 ;
      RECT 55.8 74.4 57 77.4 ;
      RECT 56.1 70.5 57 77.4 ;
      RECT 56.1 70.5 61.8 71.4 ;
      RECT 60.6 64.5 61.8 71.4 ;
      RECT 56.1 64.5 61.8 65.7 ;
      RECT 56.1 57.6 57 65.7 ;
      RECT 55.8 57.6 57 63.6 ;
      RECT 55.8 128.4 57 131.4 ;
      RECT 56.1 124.5 57 131.4 ;
      RECT 56.1 124.5 61.8 125.4 ;
      RECT 60.6 118.5 61.8 125.4 ;
      RECT 56.1 118.5 61.8 119.7 ;
      RECT 56.1 111.6 57 119.7 ;
      RECT 55.8 111.6 57 117.6 ;
      RECT 55.8 182.4 57 185.4 ;
      RECT 56.1 178.5 57 185.4 ;
      RECT 56.1 178.5 61.8 179.4 ;
      RECT 60.6 172.5 61.8 179.4 ;
      RECT 56.1 172.5 61.8 173.7 ;
      RECT 56.1 165.6 57 173.7 ;
      RECT 55.8 165.6 57 171.6 ;
      RECT 55.8 236.4 57 239.4 ;
      RECT 56.1 232.5 57 239.4 ;
      RECT 56.1 232.5 61.8 233.4 ;
      RECT 60.6 226.5 61.8 233.4 ;
      RECT 56.1 226.5 61.8 227.7 ;
      RECT 56.1 219.6 57 227.7 ;
      RECT 55.8 219.6 57 225.6 ;
      RECT 55.8 290.4 57 293.4 ;
      RECT 56.1 286.5 57 293.4 ;
      RECT 56.1 286.5 61.8 287.4 ;
      RECT 60.6 280.5 61.8 287.4 ;
      RECT 56.1 280.5 61.8 281.7 ;
      RECT 56.1 273.6 57 281.7 ;
      RECT 55.8 273.6 57 279.6 ;
      RECT 55.8 344.4 57 347.4 ;
      RECT 56.1 340.5 57 347.4 ;
      RECT 56.1 340.5 61.8 341.4 ;
      RECT 60.6 334.5 61.8 341.4 ;
      RECT 56.1 334.5 61.8 335.7 ;
      RECT 56.1 327.6 57 335.7 ;
      RECT 55.8 327.6 57 333.6 ;
      RECT 55.8 398.4 57 401.4 ;
      RECT 56.1 394.5 57 401.4 ;
      RECT 56.1 394.5 61.8 395.4 ;
      RECT 60.6 388.5 61.8 395.4 ;
      RECT 56.1 388.5 61.8 389.7 ;
      RECT 56.1 381.6 57 389.7 ;
      RECT 55.8 381.6 57 387.6 ;
      RECT 49.5 18.3 50.7 23.4 ;
      RECT 49.8 3.6 50.7 23.4 ;
      RECT 46.2 18.3 50.7 19.5 ;
      RECT 49.8 13.5 51.6 14.7 ;
      RECT 49.5 3.6 50.7 9.6 ;
      RECT 49.5 72.3 50.7 77.4 ;
      RECT 49.8 57.6 50.7 77.4 ;
      RECT 46.2 72.3 50.7 73.5 ;
      RECT 49.8 67.5 51.6 68.7 ;
      RECT 49.5 57.6 50.7 63.6 ;
      RECT 49.5 126.3 50.7 131.4 ;
      RECT 49.8 111.6 50.7 131.4 ;
      RECT 46.2 126.3 50.7 127.5 ;
      RECT 49.8 121.5 51.6 122.7 ;
      RECT 49.5 111.6 50.7 117.6 ;
      RECT 49.5 180.3 50.7 185.4 ;
      RECT 49.8 165.6 50.7 185.4 ;
      RECT 46.2 180.3 50.7 181.5 ;
      RECT 49.8 175.5 51.6 176.7 ;
      RECT 49.5 165.6 50.7 171.6 ;
      RECT 49.5 234.3 50.7 239.4 ;
      RECT 49.8 219.6 50.7 239.4 ;
      RECT 46.2 234.3 50.7 235.5 ;
      RECT 49.8 229.5 51.6 230.7 ;
      RECT 49.5 219.6 50.7 225.6 ;
      RECT 49.5 288.3 50.7 293.4 ;
      RECT 49.8 273.6 50.7 293.4 ;
      RECT 46.2 288.3 50.7 289.5 ;
      RECT 49.8 283.5 51.6 284.7 ;
      RECT 49.5 273.6 50.7 279.6 ;
      RECT 49.5 342.3 50.7 347.4 ;
      RECT 49.8 327.6 50.7 347.4 ;
      RECT 46.2 342.3 50.7 343.5 ;
      RECT 49.8 337.5 51.6 338.7 ;
      RECT 49.5 327.6 50.7 333.6 ;
      RECT 49.5 396.3 50.7 401.4 ;
      RECT 49.8 381.6 50.7 401.4 ;
      RECT 46.2 396.3 50.7 397.5 ;
      RECT 49.8 391.5 51.6 392.7 ;
      RECT 49.5 381.6 50.7 387.6 ;
      RECT 41.4 34.5 49.8 35.7 ;
      RECT 48.6 30.6 49.8 35.7 ;
      RECT 46.2 30.6 47.4 35.7 ;
      RECT 41.4 30.6 42.6 35.7 ;
      RECT 36.6 30.6 37.8 50.4 ;
      RECT 30.3 30.6 31.5 50.4 ;
      RECT 30.3 42.3 37.8 43.5 ;
      RECT 36.6 38.7 49.8 39.9 ;
      RECT 48.6 36.6 49.8 39.9 ;
      RECT 48.6 42.3 49.8 50.4 ;
      RECT 46.2 42.3 47.4 50.4 ;
      RECT 41.4 42.3 42.6 50.4 ;
      RECT 41.4 42.3 49.8 43.5 ;
      RECT 41.4 88.5 49.8 89.7 ;
      RECT 48.6 84.6 49.8 89.7 ;
      RECT 46.2 84.6 47.4 89.7 ;
      RECT 41.4 84.6 42.6 89.7 ;
      RECT 36.6 84.6 37.8 104.4 ;
      RECT 30.3 84.6 31.5 104.4 ;
      RECT 30.3 96.3 37.8 97.5 ;
      RECT 36.6 92.7 49.8 93.9 ;
      RECT 48.6 90.6 49.8 93.9 ;
      RECT 48.6 96.3 49.8 104.4 ;
      RECT 46.2 96.3 47.4 104.4 ;
      RECT 41.4 96.3 42.6 104.4 ;
      RECT 41.4 96.3 49.8 97.5 ;
      RECT 41.4 142.5 49.8 143.7 ;
      RECT 48.6 138.6 49.8 143.7 ;
      RECT 46.2 138.6 47.4 143.7 ;
      RECT 41.4 138.6 42.6 143.7 ;
      RECT 36.6 138.6 37.8 158.4 ;
      RECT 30.3 138.6 31.5 158.4 ;
      RECT 30.3 150.3 37.8 151.5 ;
      RECT 36.6 146.7 49.8 147.9 ;
      RECT 48.6 144.6 49.8 147.9 ;
      RECT 48.6 150.3 49.8 158.4 ;
      RECT 46.2 150.3 47.4 158.4 ;
      RECT 41.4 150.3 42.6 158.4 ;
      RECT 41.4 150.3 49.8 151.5 ;
      RECT 41.4 196.5 49.8 197.7 ;
      RECT 48.6 192.6 49.8 197.7 ;
      RECT 46.2 192.6 47.4 197.7 ;
      RECT 41.4 192.6 42.6 197.7 ;
      RECT 36.6 192.6 37.8 212.4 ;
      RECT 30.3 192.6 31.5 212.4 ;
      RECT 30.3 204.3 37.8 205.5 ;
      RECT 36.6 200.7 49.8 201.9 ;
      RECT 48.6 198.6 49.8 201.9 ;
      RECT 48.6 204.3 49.8 212.4 ;
      RECT 46.2 204.3 47.4 212.4 ;
      RECT 41.4 204.3 42.6 212.4 ;
      RECT 41.4 204.3 49.8 205.5 ;
      RECT 41.4 250.5 49.8 251.7 ;
      RECT 48.6 246.6 49.8 251.7 ;
      RECT 46.2 246.6 47.4 251.7 ;
      RECT 41.4 246.6 42.6 251.7 ;
      RECT 36.6 246.6 37.8 266.4 ;
      RECT 30.3 246.6 31.5 266.4 ;
      RECT 30.3 258.3 37.8 259.5 ;
      RECT 36.6 254.7 49.8 255.9 ;
      RECT 48.6 252.6 49.8 255.9 ;
      RECT 48.6 258.3 49.8 266.4 ;
      RECT 46.2 258.3 47.4 266.4 ;
      RECT 41.4 258.3 42.6 266.4 ;
      RECT 41.4 258.3 49.8 259.5 ;
      RECT 41.4 304.5 49.8 305.7 ;
      RECT 48.6 300.6 49.8 305.7 ;
      RECT 46.2 300.6 47.4 305.7 ;
      RECT 41.4 300.6 42.6 305.7 ;
      RECT 36.6 300.6 37.8 320.4 ;
      RECT 30.3 300.6 31.5 320.4 ;
      RECT 30.3 312.3 37.8 313.5 ;
      RECT 36.6 308.7 49.8 309.9 ;
      RECT 48.6 306.6 49.8 309.9 ;
      RECT 48.6 312.3 49.8 320.4 ;
      RECT 46.2 312.3 47.4 320.4 ;
      RECT 41.4 312.3 42.6 320.4 ;
      RECT 41.4 312.3 49.8 313.5 ;
      RECT 41.4 358.5 49.8 359.7 ;
      RECT 48.6 354.6 49.8 359.7 ;
      RECT 46.2 354.6 47.4 359.7 ;
      RECT 41.4 354.6 42.6 359.7 ;
      RECT 36.6 354.6 37.8 374.4 ;
      RECT 30.3 354.6 31.5 374.4 ;
      RECT 30.3 366.3 37.8 367.5 ;
      RECT 36.6 362.7 49.8 363.9 ;
      RECT 48.6 360.6 49.8 363.9 ;
      RECT 48.6 366.3 49.8 374.4 ;
      RECT 46.2 366.3 47.4 374.4 ;
      RECT 41.4 366.3 42.6 374.4 ;
      RECT 41.4 366.3 49.8 367.5 ;
      RECT 41.4 412.5 49.8 413.7 ;
      RECT 48.6 408.6 49.8 413.7 ;
      RECT 46.2 408.6 47.4 413.7 ;
      RECT 41.4 408.6 42.6 413.7 ;
      RECT 36.6 408.6 37.8 428.4 ;
      RECT 30.3 408.6 31.5 428.4 ;
      RECT 30.3 420.3 37.8 421.5 ;
      RECT 36.6 416.7 49.8 417.9 ;
      RECT 48.6 414.6 49.8 417.9 ;
      RECT 48.6 420.3 49.8 428.4 ;
      RECT 46.2 420.3 47.4 428.4 ;
      RECT 41.4 420.3 42.6 428.4 ;
      RECT 41.4 420.3 49.8 421.5 ;
      RECT 42.9 20.4 44.1 23.4 ;
      RECT 43.2 16.5 44.1 23.4 ;
      RECT 43.2 16.5 48.9 17.4 ;
      RECT 47.7 10.5 48.9 17.4 ;
      RECT 43.2 10.5 48.9 11.7 ;
      RECT 43.2 3.6 44.1 11.7 ;
      RECT 42.9 3.6 44.1 9.6 ;
      RECT 42.9 74.4 44.1 77.4 ;
      RECT 43.2 70.5 44.1 77.4 ;
      RECT 43.2 70.5 48.9 71.4 ;
      RECT 47.7 64.5 48.9 71.4 ;
      RECT 43.2 64.5 48.9 65.7 ;
      RECT 43.2 57.6 44.1 65.7 ;
      RECT 42.9 57.6 44.1 63.6 ;
      RECT 42.9 128.4 44.1 131.4 ;
      RECT 43.2 124.5 44.1 131.4 ;
      RECT 43.2 124.5 48.9 125.4 ;
      RECT 47.7 118.5 48.9 125.4 ;
      RECT 43.2 118.5 48.9 119.7 ;
      RECT 43.2 111.6 44.1 119.7 ;
      RECT 42.9 111.6 44.1 117.6 ;
      RECT 42.9 182.4 44.1 185.4 ;
      RECT 43.2 178.5 44.1 185.4 ;
      RECT 43.2 178.5 48.9 179.4 ;
      RECT 47.7 172.5 48.9 179.4 ;
      RECT 43.2 172.5 48.9 173.7 ;
      RECT 43.2 165.6 44.1 173.7 ;
      RECT 42.9 165.6 44.1 171.6 ;
      RECT 42.9 236.4 44.1 239.4 ;
      RECT 43.2 232.5 44.1 239.4 ;
      RECT 43.2 232.5 48.9 233.4 ;
      RECT 47.7 226.5 48.9 233.4 ;
      RECT 43.2 226.5 48.9 227.7 ;
      RECT 43.2 219.6 44.1 227.7 ;
      RECT 42.9 219.6 44.1 225.6 ;
      RECT 42.9 290.4 44.1 293.4 ;
      RECT 43.2 286.5 44.1 293.4 ;
      RECT 43.2 286.5 48.9 287.4 ;
      RECT 47.7 280.5 48.9 287.4 ;
      RECT 43.2 280.5 48.9 281.7 ;
      RECT 43.2 273.6 44.1 281.7 ;
      RECT 42.9 273.6 44.1 279.6 ;
      RECT 42.9 344.4 44.1 347.4 ;
      RECT 43.2 340.5 44.1 347.4 ;
      RECT 43.2 340.5 48.9 341.4 ;
      RECT 47.7 334.5 48.9 341.4 ;
      RECT 43.2 334.5 48.9 335.7 ;
      RECT 43.2 327.6 44.1 335.7 ;
      RECT 42.9 327.6 44.1 333.6 ;
      RECT 42.9 398.4 44.1 401.4 ;
      RECT 43.2 394.5 44.1 401.4 ;
      RECT 43.2 394.5 48.9 395.4 ;
      RECT 47.7 388.5 48.9 395.4 ;
      RECT 43.2 388.5 48.9 389.7 ;
      RECT 43.2 381.6 44.1 389.7 ;
      RECT 42.9 381.6 44.1 387.6 ;
      RECT 36.6 3.6 37.8 23.4 ;
      RECT 41.1 10.5 42.3 12.9 ;
      RECT 36.6 10.5 42.3 11.7 ;
      RECT 36.6 57.6 37.8 77.4 ;
      RECT 41.1 64.5 42.3 66.9 ;
      RECT 36.6 64.5 42.3 65.7 ;
      RECT 36.6 111.6 37.8 131.4 ;
      RECT 41.1 118.5 42.3 120.9 ;
      RECT 36.6 118.5 42.3 119.7 ;
      RECT 36.6 165.6 37.8 185.4 ;
      RECT 41.1 172.5 42.3 174.9 ;
      RECT 36.6 172.5 42.3 173.7 ;
      RECT 36.6 219.6 37.8 239.4 ;
      RECT 41.1 226.5 42.3 228.9 ;
      RECT 36.6 226.5 42.3 227.7 ;
      RECT 36.6 273.6 37.8 293.4 ;
      RECT 41.1 280.5 42.3 282.9 ;
      RECT 36.6 280.5 42.3 281.7 ;
      RECT 36.6 327.6 37.8 347.4 ;
      RECT 41.1 334.5 42.3 336.9 ;
      RECT 36.6 334.5 42.3 335.7 ;
      RECT 36.6 381.6 37.8 401.4 ;
      RECT 41.1 388.5 42.3 390.9 ;
      RECT 36.6 388.5 42.3 389.7 ;
      RECT 29.4 17.4 30.6 23.4 ;
      RECT 34.2 17.1 35.4 19.5 ;
      RECT 29.4 17.4 35.4 18.3 ;
      RECT 30.9 17.1 35.4 18.3 ;
      RECT 30.9 10.5 31.8 18.3 ;
      RECT 28.2 10.5 31.8 11.4 ;
      RECT 28.2 3.6 29.1 11.4 ;
      RECT 27.9 3.6 29.1 9.6 ;
      RECT 29.4 71.4 30.6 77.4 ;
      RECT 34.2 71.1 35.4 73.5 ;
      RECT 29.4 71.4 35.4 72.3 ;
      RECT 30.9 71.1 35.4 72.3 ;
      RECT 30.9 64.5 31.8 72.3 ;
      RECT 28.2 64.5 31.8 65.4 ;
      RECT 28.2 57.6 29.1 65.4 ;
      RECT 27.9 57.6 29.1 63.6 ;
      RECT 29.4 125.4 30.6 131.4 ;
      RECT 34.2 125.1 35.4 127.5 ;
      RECT 29.4 125.4 35.4 126.3 ;
      RECT 30.9 125.1 35.4 126.3 ;
      RECT 30.9 118.5 31.8 126.3 ;
      RECT 28.2 118.5 31.8 119.4 ;
      RECT 28.2 111.6 29.1 119.4 ;
      RECT 27.9 111.6 29.1 117.6 ;
      RECT 29.4 179.4 30.6 185.4 ;
      RECT 34.2 179.1 35.4 181.5 ;
      RECT 29.4 179.4 35.4 180.3 ;
      RECT 30.9 179.1 35.4 180.3 ;
      RECT 30.9 172.5 31.8 180.3 ;
      RECT 28.2 172.5 31.8 173.4 ;
      RECT 28.2 165.6 29.1 173.4 ;
      RECT 27.9 165.6 29.1 171.6 ;
      RECT 29.4 233.4 30.6 239.4 ;
      RECT 34.2 233.1 35.4 235.5 ;
      RECT 29.4 233.4 35.4 234.3 ;
      RECT 30.9 233.1 35.4 234.3 ;
      RECT 30.9 226.5 31.8 234.3 ;
      RECT 28.2 226.5 31.8 227.4 ;
      RECT 28.2 219.6 29.1 227.4 ;
      RECT 27.9 219.6 29.1 225.6 ;
      RECT 29.4 287.4 30.6 293.4 ;
      RECT 34.2 287.1 35.4 289.5 ;
      RECT 29.4 287.4 35.4 288.3 ;
      RECT 30.9 287.1 35.4 288.3 ;
      RECT 30.9 280.5 31.8 288.3 ;
      RECT 28.2 280.5 31.8 281.4 ;
      RECT 28.2 273.6 29.1 281.4 ;
      RECT 27.9 273.6 29.1 279.6 ;
      RECT 29.4 341.4 30.6 347.4 ;
      RECT 34.2 341.1 35.4 343.5 ;
      RECT 29.4 341.4 35.4 342.3 ;
      RECT 30.9 341.1 35.4 342.3 ;
      RECT 30.9 334.5 31.8 342.3 ;
      RECT 28.2 334.5 31.8 335.4 ;
      RECT 28.2 327.6 29.1 335.4 ;
      RECT 27.9 327.6 29.1 333.6 ;
      RECT 29.4 395.4 30.6 401.4 ;
      RECT 34.2 395.1 35.4 397.5 ;
      RECT 29.4 395.4 35.4 396.3 ;
      RECT 30.9 395.1 35.4 396.3 ;
      RECT 30.9 388.5 31.8 396.3 ;
      RECT 28.2 388.5 31.8 389.4 ;
      RECT 28.2 381.6 29.1 389.4 ;
      RECT 27.9 381.6 29.1 387.6 ;
      RECT 23.1 34.5 29.1 35.7 ;
      RECT 27.9 30.6 29.1 35.7 ;
      RECT 23.1 30.6 24.3 35.7 ;
      RECT 27.9 42.3 29.1 50.4 ;
      RECT 23.1 42.3 24.3 50.4 ;
      RECT 23.1 42.3 29.1 43.5 ;
      RECT 23.1 88.5 29.1 89.7 ;
      RECT 27.9 84.6 29.1 89.7 ;
      RECT 23.1 84.6 24.3 89.7 ;
      RECT 27.9 96.3 29.1 104.4 ;
      RECT 23.1 96.3 24.3 104.4 ;
      RECT 23.1 96.3 29.1 97.5 ;
      RECT 23.1 142.5 29.1 143.7 ;
      RECT 27.9 138.6 29.1 143.7 ;
      RECT 23.1 138.6 24.3 143.7 ;
      RECT 27.9 150.3 29.1 158.4 ;
      RECT 23.1 150.3 24.3 158.4 ;
      RECT 23.1 150.3 29.1 151.5 ;
      RECT 23.1 196.5 29.1 197.7 ;
      RECT 27.9 192.6 29.1 197.7 ;
      RECT 23.1 192.6 24.3 197.7 ;
      RECT 27.9 204.3 29.1 212.4 ;
      RECT 23.1 204.3 24.3 212.4 ;
      RECT 23.1 204.3 29.1 205.5 ;
      RECT 23.1 250.5 29.1 251.7 ;
      RECT 27.9 246.6 29.1 251.7 ;
      RECT 23.1 246.6 24.3 251.7 ;
      RECT 27.9 258.3 29.1 266.4 ;
      RECT 23.1 258.3 24.3 266.4 ;
      RECT 23.1 258.3 29.1 259.5 ;
      RECT 23.1 304.5 29.1 305.7 ;
      RECT 27.9 300.6 29.1 305.7 ;
      RECT 23.1 300.6 24.3 305.7 ;
      RECT 27.9 312.3 29.1 320.4 ;
      RECT 23.1 312.3 24.3 320.4 ;
      RECT 23.1 312.3 29.1 313.5 ;
      RECT 23.1 358.5 29.1 359.7 ;
      RECT 27.9 354.6 29.1 359.7 ;
      RECT 23.1 354.6 24.3 359.7 ;
      RECT 27.9 366.3 29.1 374.4 ;
      RECT 23.1 366.3 24.3 374.4 ;
      RECT 23.1 366.3 29.1 367.5 ;
      RECT 23.1 412.5 29.1 413.7 ;
      RECT 27.9 408.6 29.1 413.7 ;
      RECT 23.1 408.6 24.3 413.7 ;
      RECT 27.9 420.3 29.1 428.4 ;
      RECT 23.1 420.3 24.3 428.4 ;
      RECT 23.1 420.3 29.1 421.5 ;
      RECT 16.5 24.3 17.7 47.4 ;
      RECT 20.7 24.3 21.9 33.6 ;
      RECT 0 24.3 25.5 29.7 ;
      RECT 11.7 20.4 12.9 29.7 ;
      RECT 7.5 15.6 8.7 29.7 ;
      RECT 6.9 15.6 10.8 16.8 ;
      RECT 11.7 51.3 12.9 63.6 ;
      RECT 0 51.3 25.5 56.7 ;
      RECT 20.7 44.4 21.9 56.7 ;
      RECT 11.7 105.3 12.9 117.6 ;
      RECT 0 105.3 25.5 110.7 ;
      RECT 20.7 98.4 21.9 110.7 ;
      RECT 11.7 159.3 12.9 171.6 ;
      RECT 0 159.3 25.5 164.7 ;
      RECT 20.7 152.4 21.9 164.7 ;
      RECT 11.7 213.3 12.9 225.6 ;
      RECT 0 213.3 25.5 218.7 ;
      RECT 20.7 206.4 21.9 218.7 ;
      RECT 11.7 267.3 12.9 279.6 ;
      RECT 0 267.3 25.5 272.7 ;
      RECT 20.7 260.4 21.9 272.7 ;
      RECT 11.7 321.3 12.9 333.6 ;
      RECT 0 321.3 25.5 326.7 ;
      RECT 20.7 314.4 21.9 326.7 ;
      RECT 11.7 375.3 12.9 387.6 ;
      RECT 0 375.3 25.5 380.7 ;
      RECT 20.7 368.4 21.9 380.7 ;
      RECT 16.5 402.3 17.7 425.4 ;
      RECT 20.7 402.3 21.9 411.6 ;
      RECT 0 402.3 25.5 407.7 ;
      RECT 11.7 398.4 12.9 407.7 ;
      RECT 7.5 393.6 8.7 407.7 ;
      RECT 6.9 393.6 10.8 394.8 ;
      RECT 7.8 429.3 25.5 430.2 ;
      RECT 20.7 422.4 21.9 430.2 ;
      RECT 11.7 30.6 12.9 47.4 ;
      RECT 6.9 30.6 12.9 31.8 ;
      RECT 11.7 84.6 12.9 101.4 ;
      RECT 6.9 84.6 12.9 85.8 ;
      RECT 11.7 138.6 12.9 155.4 ;
      RECT 6.9 138.6 12.9 139.8 ;
      RECT 11.7 192.6 12.9 209.4 ;
      RECT 6.9 192.6 12.9 193.8 ;
      RECT 11.7 246.6 12.9 263.4 ;
      RECT 6.9 246.6 12.9 247.8 ;
      RECT 11.7 300.6 12.9 317.4 ;
      RECT 6.9 300.6 12.9 301.8 ;
      RECT 11.7 354.6 12.9 371.4 ;
      RECT 6.9 354.6 12.9 355.8 ;
      RECT 11.7 408.6 12.9 425.4 ;
      RECT 6.9 408.6 12.9 409.8 ;
      RECT 139.2 3.6 140.7 9.6 ;
      RECT 135.9 13.2 137.1 15.6 ;
      RECT 135.9 67.2 137.1 69.6 ;
      RECT 135.9 121.2 137.1 123.6 ;
      RECT 135.9 175.2 137.1 177.6 ;
      RECT 135.9 229.2 137.1 231.6 ;
      RECT 135.9 283.2 137.1 285.6 ;
      RECT 135.9 337.2 137.1 339.6 ;
      RECT 135.9 391.2 137.1 393.6 ;
      RECT 132.3 13.5 134.7 14.7 ;
      RECT 132.3 67.5 134.7 68.7 ;
      RECT 132.3 121.5 134.7 122.7 ;
      RECT 132.3 175.5 134.7 176.7 ;
      RECT 132.3 229.5 134.7 230.7 ;
      RECT 132.3 283.5 134.7 284.7 ;
      RECT 132.3 337.5 134.7 338.7 ;
      RECT 132.3 391.5 134.7 392.7 ;
      RECT 131.7 15.9 132.9 18.3 ;
      RECT 131.7 69.9 132.9 72.3 ;
      RECT 131.7 123.9 132.9 126.3 ;
      RECT 131.7 177.9 132.9 180.3 ;
      RECT 131.7 231.9 132.9 234.3 ;
      RECT 131.7 285.9 132.9 288.3 ;
      RECT 131.7 339.9 132.9 342.3 ;
      RECT 131.7 393.9 132.9 396.3 ;
      RECT 131.4 3.6 132.6 9.6 ;
      RECT 126.3 3.6 127.8 9.6 ;
      RECT 123 13.2 124.2 15.6 ;
      RECT 123 67.2 124.2 69.6 ;
      RECT 123 121.2 124.2 123.6 ;
      RECT 123 175.2 124.2 177.6 ;
      RECT 123 229.2 124.2 231.6 ;
      RECT 123 283.2 124.2 285.6 ;
      RECT 123 337.2 124.2 339.6 ;
      RECT 123 391.2 124.2 393.6 ;
      RECT 118.8 17.1 120 19.5 ;
      RECT 118.8 71.1 120 73.5 ;
      RECT 118.8 125.1 120 127.5 ;
      RECT 118.8 179.1 120 181.5 ;
      RECT 118.8 233.1 120 235.5 ;
      RECT 118.8 287.1 120 289.5 ;
      RECT 118.8 341.1 120 343.5 ;
      RECT 118.8 395.1 120 397.5 ;
      RECT 118.5 3.6 119.7 9.6 ;
      RECT 118.2 13.5 119.4 15.9 ;
      RECT 118.2 67.5 119.4 69.9 ;
      RECT 118.2 121.5 119.4 123.9 ;
      RECT 118.2 175.5 119.4 177.9 ;
      RECT 118.2 229.5 119.4 231.9 ;
      RECT 118.2 283.5 119.4 285.9 ;
      RECT 118.2 337.5 119.4 339.9 ;
      RECT 118.2 391.5 119.4 393.9 ;
      RECT 112.2 3.6 113.4 9.6 ;
      RECT 111.9 31.2 113.1 44.4 ;
      RECT 111.9 85.2 113.1 98.4 ;
      RECT 111.9 139.2 113.1 152.4 ;
      RECT 111.9 193.2 113.1 206.4 ;
      RECT 111.9 247.2 113.1 260.4 ;
      RECT 111.9 301.2 113.1 314.4 ;
      RECT 111.9 355.2 113.1 368.4 ;
      RECT 111.9 409.2 113.1 422.4 ;
      RECT 109.8 3.6 111 9.6 ;
      RECT 109.8 33.6 111 47.4 ;
      RECT 109.8 87.6 111 101.4 ;
      RECT 109.8 141.6 111 155.4 ;
      RECT 109.8 195.6 111 209.4 ;
      RECT 109.8 249.6 111 263.4 ;
      RECT 109.8 303.6 111 317.4 ;
      RECT 109.8 357.6 111 371.4 ;
      RECT 109.8 411.6 111 425.4 ;
      RECT 105 12.3 109.5 13.5 ;
      RECT 105 66.3 109.5 67.5 ;
      RECT 105 120.3 109.5 121.5 ;
      RECT 105 174.3 109.5 175.5 ;
      RECT 105 228.3 109.5 229.5 ;
      RECT 105 282.3 109.5 283.5 ;
      RECT 105 336.3 109.5 337.5 ;
      RECT 105 390.3 109.5 391.5 ;
      RECT 107.4 32.4 108.6 47.4 ;
      RECT 107.4 86.4 108.6 101.4 ;
      RECT 107.4 140.4 108.6 155.4 ;
      RECT 107.4 194.4 108.6 209.4 ;
      RECT 107.4 248.4 108.6 263.4 ;
      RECT 107.4 302.4 108.6 317.4 ;
      RECT 107.4 356.4 108.6 371.4 ;
      RECT 107.4 410.4 108.6 425.4 ;
      RECT 105.6 15.3 108.3 16.5 ;
      RECT 105.6 69.3 108.3 70.5 ;
      RECT 105.6 123.3 108.3 124.5 ;
      RECT 105.6 177.3 108.3 178.5 ;
      RECT 105.6 231.3 108.3 232.5 ;
      RECT 105.6 285.3 108.3 286.5 ;
      RECT 105.6 339.3 108.3 340.5 ;
      RECT 105.6 393.3 108.3 394.5 ;
      RECT 105.3 48.9 107.7 50.1 ;
      RECT 105.3 102.9 107.7 104.1 ;
      RECT 105.3 156.9 107.7 158.1 ;
      RECT 105.3 210.9 107.7 212.1 ;
      RECT 105.3 264.9 107.7 266.1 ;
      RECT 105.3 318.9 107.7 320.1 ;
      RECT 105.3 372.9 107.7 374.1 ;
      RECT 105.3 426.9 107.7 428.1 ;
      RECT 105 3.6 106.2 9.6 ;
      RECT 102.9 9.6 104.1 22.8 ;
      RECT 102.9 63.6 104.1 76.8 ;
      RECT 102.9 117.6 104.1 130.8 ;
      RECT 102.9 171.6 104.1 184.8 ;
      RECT 102.9 225.6 104.1 238.8 ;
      RECT 102.9 279.6 104.1 292.8 ;
      RECT 102.9 333.6 104.1 346.8 ;
      RECT 102.9 387.6 104.1 400.8 ;
      RECT 102.6 30.6 103.8 50.4 ;
      RECT 102.6 84.6 103.8 104.4 ;
      RECT 102.6 138.6 103.8 158.4 ;
      RECT 102.6 192.6 103.8 212.4 ;
      RECT 102.6 246.6 103.8 266.4 ;
      RECT 102.6 300.6 103.8 320.4 ;
      RECT 102.6 354.6 103.8 374.4 ;
      RECT 102.6 408.6 103.8 428.4 ;
      RECT 100.8 6.6 102 20.4 ;
      RECT 100.8 60.6 102 74.4 ;
      RECT 100.8 114.6 102 128.4 ;
      RECT 100.8 168.6 102 182.4 ;
      RECT 100.8 222.6 102 236.4 ;
      RECT 100.8 276.6 102 290.4 ;
      RECT 100.8 330.6 102 344.4 ;
      RECT 100.8 384.6 102 398.4 ;
      RECT 100.5 40.2 101.7 42.6 ;
      RECT 100.5 94.2 101.7 96.6 ;
      RECT 100.5 148.2 101.7 150.6 ;
      RECT 100.5 202.2 101.7 204.6 ;
      RECT 100.5 256.2 101.7 258.6 ;
      RECT 100.5 310.2 101.7 312.6 ;
      RECT 100.5 364.2 101.7 366.6 ;
      RECT 100.5 418.2 101.7 420.6 ;
      RECT 100.2 422.4 101.4 428.4 ;
      RECT 98.4 6.6 99.6 23.4 ;
      RECT 98.4 60.6 99.6 77.4 ;
      RECT 98.4 114.6 99.6 131.4 ;
      RECT 98.4 168.6 99.6 185.4 ;
      RECT 98.4 222.6 99.6 239.4 ;
      RECT 98.4 276.6 99.6 293.4 ;
      RECT 98.4 330.6 99.6 347.4 ;
      RECT 98.4 384.6 99.6 401.4 ;
      RECT 98.1 30.6 99.3 44.4 ;
      RECT 98.1 84.6 99.3 98.4 ;
      RECT 98.1 138.6 99.3 152.4 ;
      RECT 98.1 192.6 99.3 206.4 ;
      RECT 98.1 246.6 99.3 260.4 ;
      RECT 98.1 300.6 99.3 314.4 ;
      RECT 98.1 354.6 99.3 368.4 ;
      RECT 98.1 408.6 99.3 422.4 ;
      RECT 96.3 3.9 98.7 5.1 ;
      RECT 96.3 57.9 98.7 59.1 ;
      RECT 96.3 111.9 98.7 113.1 ;
      RECT 96.3 165.9 98.7 167.1 ;
      RECT 96.3 219.9 98.7 221.1 ;
      RECT 96.3 273.9 98.7 275.1 ;
      RECT 96.3 327.9 98.7 329.1 ;
      RECT 96.3 381.9 98.7 383.1 ;
      RECT 87.3 429.3 98.1 430.2 ;
      RECT 96 6.6 97.2 20.4 ;
      RECT 96 33.6 97.2 47.4 ;
      RECT 96 60.6 97.2 74.4 ;
      RECT 96 87.6 97.2 101.4 ;
      RECT 96 114.6 97.2 128.4 ;
      RECT 96 141.6 97.2 155.4 ;
      RECT 96 168.6 97.2 182.4 ;
      RECT 96 195.6 97.2 209.4 ;
      RECT 96 222.6 97.2 236.4 ;
      RECT 96 249.6 97.2 263.4 ;
      RECT 96 276.6 97.2 290.4 ;
      RECT 96 303.6 97.2 317.4 ;
      RECT 96 330.6 97.2 344.4 ;
      RECT 96 357.6 97.2 371.4 ;
      RECT 96 384.6 97.2 398.4 ;
      RECT 96 411.6 97.2 425.4 ;
      RECT 93.6 3.6 94.8 23.4 ;
      RECT 93.6 32.4 94.8 47.4 ;
      RECT 93.6 57.6 94.8 77.4 ;
      RECT 93.6 86.4 94.8 101.4 ;
      RECT 93.6 111.6 94.8 131.4 ;
      RECT 93.6 140.4 94.8 155.4 ;
      RECT 93.6 165.6 94.8 185.4 ;
      RECT 93.6 194.4 94.8 209.4 ;
      RECT 93.6 219.6 94.8 239.4 ;
      RECT 93.6 248.4 94.8 263.4 ;
      RECT 93.6 273.6 94.8 293.4 ;
      RECT 93.6 302.4 94.8 317.4 ;
      RECT 93.6 327.6 94.8 347.4 ;
      RECT 93.6 356.4 94.8 371.4 ;
      RECT 93.6 381.6 94.8 401.4 ;
      RECT 93.6 410.4 94.8 425.4 ;
      RECT 86.4 48.9 93.9 50.1 ;
      RECT 86.4 102.9 93.9 104.1 ;
      RECT 86.4 156.9 93.9 158.1 ;
      RECT 86.4 210.9 93.9 212.1 ;
      RECT 86.4 264.9 93.9 266.1 ;
      RECT 86.4 318.9 93.9 320.1 ;
      RECT 86.4 372.9 93.9 374.1 ;
      RECT 86.4 426.9 93.9 428.1 ;
      RECT 91.2 3.6 92.4 9.6 ;
      RECT 89.1 18.3 92.4 19.5 ;
      RECT 89.1 72.3 92.4 73.5 ;
      RECT 89.1 126.3 92.4 127.5 ;
      RECT 89.1 180.3 92.4 181.5 ;
      RECT 89.1 234.3 92.4 235.5 ;
      RECT 89.1 288.3 92.4 289.5 ;
      RECT 89.1 342.3 92.4 343.5 ;
      RECT 89.1 396.3 92.4 397.5 ;
      RECT 78.6 6 90.3 7.2 ;
      RECT 80.7 8.1 90.3 9.3 ;
      RECT 84.9 13.5 90.3 14.7 ;
      RECT 84.9 15.6 90.3 16.8 ;
      RECT 82.8 41.4 90.3 42.6 ;
      RECT 78.6 60 90.3 61.2 ;
      RECT 80.7 62.1 90.3 63.3 ;
      RECT 84.9 67.5 90.3 68.7 ;
      RECT 84.9 69.6 90.3 70.8 ;
      RECT 82.8 95.4 90.3 96.6 ;
      RECT 78.6 114 90.3 115.2 ;
      RECT 80.7 116.1 90.3 117.3 ;
      RECT 84.9 121.5 90.3 122.7 ;
      RECT 84.9 123.6 90.3 124.8 ;
      RECT 82.8 149.4 90.3 150.6 ;
      RECT 78.6 168 90.3 169.2 ;
      RECT 80.7 170.1 90.3 171.3 ;
      RECT 84.9 175.5 90.3 176.7 ;
      RECT 84.9 177.6 90.3 178.8 ;
      RECT 82.8 203.4 90.3 204.6 ;
      RECT 78.6 222 90.3 223.2 ;
      RECT 80.7 224.1 90.3 225.3 ;
      RECT 84.9 229.5 90.3 230.7 ;
      RECT 84.9 231.6 90.3 232.8 ;
      RECT 82.8 257.4 90.3 258.6 ;
      RECT 78.6 276 90.3 277.2 ;
      RECT 80.7 278.1 90.3 279.3 ;
      RECT 84.9 283.5 90.3 284.7 ;
      RECT 84.9 285.6 90.3 286.8 ;
      RECT 82.8 311.4 90.3 312.6 ;
      RECT 78.6 330 90.3 331.2 ;
      RECT 80.7 332.1 90.3 333.3 ;
      RECT 84.9 337.5 90.3 338.7 ;
      RECT 84.9 339.6 90.3 340.8 ;
      RECT 82.8 365.4 90.3 366.6 ;
      RECT 78.6 384 90.3 385.2 ;
      RECT 80.7 386.1 90.3 387.3 ;
      RECT 84.9 391.5 90.3 392.7 ;
      RECT 84.9 393.6 90.3 394.8 ;
      RECT 66 30.6 67.2 33.6 ;
      RECT 66 35.4 67.2 37.8 ;
      RECT 66 89.4 67.2 91.8 ;
      RECT 66 143.4 67.2 145.8 ;
      RECT 66 197.4 67.2 199.8 ;
      RECT 66 251.4 67.2 253.8 ;
      RECT 66 305.4 67.2 307.8 ;
      RECT 66 359.4 67.2 361.8 ;
      RECT 66 408.6 67.2 411.6 ;
      RECT 66 413.4 67.2 415.8 ;
      RECT 63.9 3.6 65.1 17.4 ;
      RECT 63.9 20.4 65.1 23.4 ;
      RECT 63.9 57.6 65.1 71.4 ;
      RECT 63.9 74.4 65.1 77.4 ;
      RECT 63.9 111.6 65.1 125.4 ;
      RECT 63.9 128.4 65.1 131.4 ;
      RECT 63.9 165.6 65.1 179.4 ;
      RECT 63.9 182.4 65.1 185.4 ;
      RECT 63.9 219.6 65.1 233.4 ;
      RECT 63.9 236.4 65.1 239.4 ;
      RECT 63.9 273.6 65.1 287.4 ;
      RECT 63.9 290.4 65.1 293.4 ;
      RECT 63.9 327.6 65.1 341.4 ;
      RECT 63.9 344.4 65.1 347.4 ;
      RECT 63.9 381.6 65.1 395.4 ;
      RECT 63.9 398.4 65.1 401.4 ;
      RECT 63.6 30.6 64.8 50.4 ;
      RECT 63.6 84.6 64.8 104.4 ;
      RECT 63.6 138.6 64.8 158.4 ;
      RECT 63.6 192.6 64.8 212.4 ;
      RECT 63.6 246.6 64.8 266.4 ;
      RECT 63.6 300.6 64.8 320.4 ;
      RECT 63.6 354.6 64.8 374.4 ;
      RECT 63.6 408.6 64.8 428.4 ;
      RECT 59.1 18.3 63 19.5 ;
      RECT 59.1 72.3 63 73.5 ;
      RECT 59.1 126.3 63 127.5 ;
      RECT 59.1 180.3 63 181.5 ;
      RECT 59.1 234.3 63 235.5 ;
      RECT 59.1 288.3 63 289.5 ;
      RECT 59.1 342.3 63 343.5 ;
      RECT 59.1 396.3 63 397.5 ;
      RECT 61.2 30.6 62.4 33.6 ;
      RECT 61.2 408.6 62.4 411.6 ;
      RECT 59.7 3.6 61.2 9.6 ;
      RECT 59.7 20.4 61.2 23.4 ;
      RECT 59.7 398.4 61.2 401.4 ;
      RECT 55.5 37.5 57.9 38.7 ;
      RECT 55.5 91.5 57.9 92.7 ;
      RECT 55.5 145.5 57.9 146.7 ;
      RECT 55.5 199.5 57.9 200.7 ;
      RECT 55.5 253.5 57.9 254.7 ;
      RECT 55.5 307.5 57.9 308.7 ;
      RECT 55.5 361.5 57.9 362.7 ;
      RECT 55.5 415.5 57.9 416.7 ;
      RECT 56.4 13.2 57.6 15.6 ;
      RECT 56.4 67.2 57.6 69.6 ;
      RECT 56.4 121.2 57.6 123.6 ;
      RECT 56.4 175.2 57.6 177.6 ;
      RECT 56.4 229.2 57.6 231.6 ;
      RECT 56.4 283.2 57.6 285.6 ;
      RECT 56.4 337.2 57.6 339.6 ;
      RECT 56.4 391.2 57.6 393.6 ;
      RECT 54 39.9 56.4 41.1 ;
      RECT 54 93.9 56.4 95.1 ;
      RECT 54 147.9 56.4 149.1 ;
      RECT 54 201.9 56.4 203.1 ;
      RECT 54 255.9 56.4 257.1 ;
      RECT 54 309.9 56.4 311.1 ;
      RECT 54 363.9 56.4 365.1 ;
      RECT 54 417.9 56.4 419.1 ;
      RECT 52.8 13.5 55.2 14.7 ;
      RECT 52.8 42.3 55.2 43.5 ;
      RECT 52.8 67.5 55.2 68.7 ;
      RECT 52.8 96.3 55.2 97.5 ;
      RECT 52.8 121.5 55.2 122.7 ;
      RECT 52.8 150.3 55.2 151.5 ;
      RECT 52.8 175.5 55.2 176.7 ;
      RECT 52.8 204.3 55.2 205.5 ;
      RECT 52.8 229.5 55.2 230.7 ;
      RECT 52.8 258.3 55.2 259.5 ;
      RECT 52.8 283.5 55.2 284.7 ;
      RECT 52.8 312.3 55.2 313.5 ;
      RECT 52.8 337.5 55.2 338.7 ;
      RECT 52.8 366.3 55.2 367.5 ;
      RECT 52.8 391.5 55.2 392.7 ;
      RECT 52.8 420.3 55.2 421.5 ;
      RECT 53.4 30.6 54.6 33.6 ;
      RECT 53.4 408.6 54.6 411.6 ;
      RECT 52.2 15.9 53.4 18.3 ;
      RECT 52.2 69.9 53.4 72.3 ;
      RECT 52.2 123.9 53.4 126.3 ;
      RECT 52.2 177.9 53.4 180.3 ;
      RECT 52.2 231.9 53.4 234.3 ;
      RECT 52.2 285.9 53.4 288.3 ;
      RECT 52.2 339.9 53.4 342.3 ;
      RECT 52.2 393.9 53.4 396.3 ;
      RECT 51.9 3.6 53.1 9.6 ;
      RECT 51.9 20.4 53.1 23.4 ;
      RECT 51.9 398.4 53.1 401.4 ;
      RECT 46.8 3.6 48.3 9.6 ;
      RECT 46.8 20.4 48.3 23.4 ;
      RECT 46.8 398.4 48.3 401.4 ;
      RECT 44.4 36.6 46.8 37.8 ;
      RECT 44.4 90.6 46.8 91.8 ;
      RECT 44.4 144.6 46.8 145.8 ;
      RECT 44.4 198.6 46.8 199.8 ;
      RECT 44.4 252.6 46.8 253.8 ;
      RECT 44.4 306.6 46.8 307.8 ;
      RECT 44.4 360.6 46.8 361.8 ;
      RECT 44.4 414.6 46.8 415.8 ;
      RECT 43.8 30.6 45 33.6 ;
      RECT 43.8 408.6 45 411.6 ;
      RECT 43.5 13.2 44.7 15.6 ;
      RECT 43.5 67.2 44.7 69.6 ;
      RECT 43.5 121.2 44.7 123.6 ;
      RECT 43.5 175.2 44.7 177.6 ;
      RECT 43.5 229.2 44.7 231.6 ;
      RECT 43.5 283.2 44.7 285.6 ;
      RECT 43.5 337.2 44.7 339.6 ;
      RECT 43.5 391.2 44.7 393.6 ;
      RECT 39 36.6 43.5 37.8 ;
      RECT 39 90.6 43.5 91.8 ;
      RECT 39 144.6 43.5 145.8 ;
      RECT 39 198.6 43.5 199.8 ;
      RECT 39 252.6 43.5 253.8 ;
      RECT 39 306.6 43.5 307.8 ;
      RECT 39 360.6 43.5 361.8 ;
      RECT 39 414.6 43.5 415.8 ;
      RECT 39.3 17.1 40.5 19.5 ;
      RECT 39.3 71.1 40.5 73.5 ;
      RECT 39.3 125.1 40.5 127.5 ;
      RECT 39.3 179.1 40.5 181.5 ;
      RECT 39.3 233.1 40.5 235.5 ;
      RECT 39.3 287.1 40.5 289.5 ;
      RECT 39.3 341.1 40.5 343.5 ;
      RECT 39.3 395.1 40.5 397.5 ;
      RECT 39 3.6 40.2 9.6 ;
      RECT 39 20.4 40.2 23.4 ;
      RECT 39 30.6 40.2 33.6 ;
      RECT 39 41.1 40.2 43.5 ;
      RECT 39 95.1 40.2 97.5 ;
      RECT 39 149.1 40.2 151.5 ;
      RECT 39 203.1 40.2 205.5 ;
      RECT 39 257.1 40.2 259.5 ;
      RECT 39 311.1 40.2 313.5 ;
      RECT 39 365.1 40.2 367.5 ;
      RECT 39 398.4 40.2 401.4 ;
      RECT 39 408.6 40.2 411.6 ;
      RECT 39 419.1 40.2 421.5 ;
      RECT 38.7 13.5 39.9 15.9 ;
      RECT 38.7 67.5 39.9 69.9 ;
      RECT 38.7 121.5 39.9 123.9 ;
      RECT 38.7 175.5 39.9 177.9 ;
      RECT 38.7 229.5 39.9 231.9 ;
      RECT 38.7 283.5 39.9 285.9 ;
      RECT 38.7 337.5 39.9 339.9 ;
      RECT 38.7 391.5 39.9 393.9 ;
      RECT 34.5 34.5 35.7 36.9 ;
      RECT 34.5 88.5 35.7 90.9 ;
      RECT 34.5 142.5 35.7 144.9 ;
      RECT 34.5 196.5 35.7 198.9 ;
      RECT 34.5 250.5 35.7 252.9 ;
      RECT 34.5 304.5 35.7 306.9 ;
      RECT 34.5 358.5 35.7 360.9 ;
      RECT 34.5 412.5 35.7 414.9 ;
      RECT 32.7 3.6 33.9 9.6 ;
      RECT 32.7 20.4 33.9 23.4 ;
      RECT 32.7 30.6 33.9 33.6 ;
      RECT 32.7 38.7 33.9 41.1 ;
      RECT 32.7 92.7 33.9 95.1 ;
      RECT 32.7 146.7 33.9 149.1 ;
      RECT 32.7 200.7 33.9 203.1 ;
      RECT 32.7 254.7 33.9 257.1 ;
      RECT 32.7 308.7 33.9 311.1 ;
      RECT 32.7 362.7 33.9 365.1 ;
      RECT 32.7 398.4 33.9 401.4 ;
      RECT 32.7 408.6 33.9 411.6 ;
      RECT 32.7 416.7 33.9 419.1 ;
      RECT 30.3 3.6 31.5 9.6 ;
      RECT 25.5 12.3 30 13.5 ;
      RECT 25.5 66.3 30 67.5 ;
      RECT 25.5 120.3 30 121.5 ;
      RECT 25.5 174.3 30 175.5 ;
      RECT 25.5 228.3 30 229.5 ;
      RECT 25.5 282.3 30 283.5 ;
      RECT 25.5 336.3 30 337.5 ;
      RECT 25.5 390.3 30 391.5 ;
      RECT 26.7 40.2 29.1 41.4 ;
      RECT 26.7 94.2 29.1 95.4 ;
      RECT 26.7 148.2 29.1 149.4 ;
      RECT 26.7 202.2 29.1 203.4 ;
      RECT 26.7 256.2 29.1 257.4 ;
      RECT 26.7 310.2 29.1 311.4 ;
      RECT 26.7 364.2 29.1 365.4 ;
      RECT 26.7 418.2 29.1 419.4 ;
      RECT 26.1 15.3 28.8 16.5 ;
      RECT 26.1 69.3 28.8 70.5 ;
      RECT 26.1 123.3 28.8 124.5 ;
      RECT 26.1 177.3 28.8 178.5 ;
      RECT 26.1 231.3 28.8 232.5 ;
      RECT 26.1 285.3 28.8 286.5 ;
      RECT 26.1 339.3 28.8 340.5 ;
      RECT 26.1 393.3 28.8 394.5 ;
      RECT 25.5 36.6 27.9 37.8 ;
      RECT 25.5 90.6 27.9 91.8 ;
      RECT 25.5 144.6 27.9 145.8 ;
      RECT 25.5 198.6 27.9 199.8 ;
      RECT 25.5 252.6 27.9 253.8 ;
      RECT 25.5 306.6 27.9 307.8 ;
      RECT 25.5 360.6 27.9 361.8 ;
      RECT 25.5 414.6 27.9 415.8 ;
      RECT 25.5 3.6 26.7 9.6 ;
      RECT 25.5 17.4 26.7 23.4 ;
      RECT 25.5 30.6 26.7 33.6 ;
      RECT 25.5 44.4 26.7 50.4 ;
      RECT 25.5 57.6 26.7 63.6 ;
      RECT 25.5 98.4 26.7 104.4 ;
      RECT 25.5 111.6 26.7 117.6 ;
      RECT 25.5 152.4 26.7 158.4 ;
      RECT 25.5 165.6 26.7 171.6 ;
      RECT 25.5 206.4 26.7 212.4 ;
      RECT 25.5 219.6 26.7 225.6 ;
      RECT 25.5 260.4 26.7 266.4 ;
      RECT 25.5 273.6 26.7 279.6 ;
      RECT 25.5 314.4 26.7 320.4 ;
      RECT 25.5 327.6 26.7 333.6 ;
      RECT 25.5 368.4 26.7 374.4 ;
      RECT 25.5 381.6 26.7 387.6 ;
      RECT 25.5 395.4 26.7 401.4 ;
      RECT 25.5 408.6 26.7 411.6 ;
      RECT 25.5 422.4 26.7 428.4 ;
      RECT 23.4 9.6 24.6 22.8 ;
      RECT 23.4 63.6 24.6 76.8 ;
      RECT 23.4 117.6 24.6 130.8 ;
      RECT 23.4 171.6 24.6 184.8 ;
      RECT 23.4 225.6 24.6 238.8 ;
      RECT 23.4 279.6 24.6 292.8 ;
      RECT 23.4 333.6 24.6 346.8 ;
      RECT 23.4 387.6 24.6 400.8 ;
      RECT 21.3 6.6 22.5 20.4 ;
      RECT 21.3 60.6 22.5 74.4 ;
      RECT 21.3 114.6 22.5 128.4 ;
      RECT 21.3 168.6 22.5 182.4 ;
      RECT 21.3 222.6 22.5 236.4 ;
      RECT 21.3 276.6 22.5 290.4 ;
      RECT 21.3 330.6 22.5 344.4 ;
      RECT 21.3 384.6 22.5 398.4 ;
      RECT 20.7 34.5 21.9 36.9 ;
      RECT 20.7 88.5 21.9 90.9 ;
      RECT 20.7 142.5 21.9 144.9 ;
      RECT 20.7 196.5 21.9 198.9 ;
      RECT 20.7 250.5 21.9 252.9 ;
      RECT 20.7 304.5 21.9 306.9 ;
      RECT 20.7 358.5 21.9 360.9 ;
      RECT 20.7 412.5 21.9 414.9 ;
      RECT 18.9 6.6 20.1 23.4 ;
      RECT 18.9 60.6 20.1 77.4 ;
      RECT 18.9 114.6 20.1 131.4 ;
      RECT 18.9 168.6 20.1 185.4 ;
      RECT 18.9 222.6 20.1 239.4 ;
      RECT 18.9 276.6 20.1 293.4 ;
      RECT 18.9 330.6 20.1 347.4 ;
      RECT 18.9 384.6 20.1 401.4 ;
      RECT 18.6 30.6 19.8 44.4 ;
      RECT 18.6 84.6 19.8 98.4 ;
      RECT 18.6 138.6 19.8 152.4 ;
      RECT 18.6 192.6 19.8 206.4 ;
      RECT 18.6 246.6 19.8 260.4 ;
      RECT 18.6 300.6 19.8 314.4 ;
      RECT 18.6 354.6 19.8 368.4 ;
      RECT 18.6 408.6 19.8 422.4 ;
      RECT 16.8 3.9 19.2 5.1 ;
      RECT 16.8 57.9 19.2 59.1 ;
      RECT 16.8 111.9 19.2 113.1 ;
      RECT 16.8 165.9 19.2 167.1 ;
      RECT 16.8 219.9 19.2 221.1 ;
      RECT 16.8 273.9 19.2 275.1 ;
      RECT 16.8 327.9 19.2 329.1 ;
      RECT 16.8 381.9 19.2 383.1 ;
      RECT 16.5 6.6 17.7 20.4 ;
      RECT 16.5 60.6 17.7 74.4 ;
      RECT 16.5 114.6 17.7 128.4 ;
      RECT 16.5 168.6 17.7 182.4 ;
      RECT 16.5 222.6 17.7 236.4 ;
      RECT 16.5 276.6 17.7 290.4 ;
      RECT 16.5 330.6 17.7 344.4 ;
      RECT 16.5 384.6 17.7 398.4 ;
      RECT 14.1 3.6 15.3 23.4 ;
      RECT 14.1 33.6 15.3 47.4 ;
      RECT 14.1 57.6 15.3 77.4 ;
      RECT 14.1 87.6 15.3 101.4 ;
      RECT 14.1 111.6 15.3 131.4 ;
      RECT 14.1 141.6 15.3 155.4 ;
      RECT 14.1 165.6 15.3 185.4 ;
      RECT 14.1 195.6 15.3 209.4 ;
      RECT 14.1 219.6 15.3 239.4 ;
      RECT 14.1 249.6 15.3 263.4 ;
      RECT 14.1 273.6 15.3 293.4 ;
      RECT 14.1 303.6 15.3 317.4 ;
      RECT 14.1 327.6 15.3 347.4 ;
      RECT 14.1 357.6 15.3 371.4 ;
      RECT 14.1 381.6 15.3 401.4 ;
      RECT 14.1 411.6 15.3 425.4 ;
      RECT 6.9 48.9 14.4 50.1 ;
      RECT 6.9 102.9 14.4 104.1 ;
      RECT 6.9 156.9 14.4 158.1 ;
      RECT 6.9 210.9 14.4 212.1 ;
      RECT 6.9 264.9 14.4 266.1 ;
      RECT 6.9 318.9 14.4 320.1 ;
      RECT 6.9 372.9 14.4 374.1 ;
      RECT 6.9 426.9 14.4 428.1 ;
      RECT 11.7 3.6 12.9 9.6 ;
      RECT 9.6 18.3 12.9 19.5 ;
      RECT 9.6 72.3 12.9 73.5 ;
      RECT 9.6 126.3 12.9 127.5 ;
      RECT 9.6 180.3 12.9 181.5 ;
      RECT 9.6 234.3 12.9 235.5 ;
      RECT 9.6 288.3 12.9 289.5 ;
      RECT 9.6 342.3 12.9 343.5 ;
      RECT 9.6 396.3 12.9 397.5 ;
      RECT 0.9 6 10.8 7.2 ;
      RECT 3 8.1 10.8 9.3 ;
      RECT 5.4 13.5 10.8 14.7 ;
      RECT 0.9 60 10.8 61.2 ;
      RECT 3 62.1 10.8 63.3 ;
      RECT 5.4 67.5 10.8 68.7 ;
      RECT 0.9 114 10.8 115.2 ;
      RECT 3 116.1 10.8 117.3 ;
      RECT 5.4 121.5 10.8 122.7 ;
      RECT 0.9 168 10.8 169.2 ;
      RECT 3 170.1 10.8 171.3 ;
      RECT 5.4 175.5 10.8 176.7 ;
      RECT 0.9 222 10.8 223.2 ;
      RECT 3 224.1 10.8 225.3 ;
      RECT 5.4 229.5 10.8 230.7 ;
      RECT 0.9 276 10.8 277.2 ;
      RECT 3 278.1 10.8 279.3 ;
      RECT 5.4 283.5 10.8 284.7 ;
      RECT 0.9 330 10.8 331.2 ;
      RECT 3 332.1 10.8 333.3 ;
      RECT 5.4 337.5 10.8 338.7 ;
      RECT 0.9 384 10.8 385.2 ;
      RECT 3 386.1 10.8 387.3 ;
      RECT 5.4 391.5 10.8 392.7 ;
  END
END bpm_custom

END LIBRARY
