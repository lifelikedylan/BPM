* SPICE NETLIST
***************************************

.SUBCKT ______inv_magic_inverter A gnd vdd Y
** N=4 EP=4 IP=0 FDC=2
M0 Y A gnd gnd n L=6e-07 W=3e-06 AD=4.5e-12 AS=4.5e-12 PD=9e-06 PS=9e-06 $X=2100 $Y=2400 $D=1
M1 Y A vdd vdd p L=6e-07 W=6e-06 AD=9e-12 AS=9e-12 PD=1.5e-05 PS=1.5e-05 $X=2100 $Y=16200 $D=0
.ENDS
***************************************
.SUBCKT bs1 en clk fa_in Cout Out Cin
** N=48 EP=6 IP=8 FDC=70
M0 11 8 5 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=12600 $Y=16500 $D=1
M1 12 9 6 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=12600 $Y=32700 $D=1
M2 3 4 11 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=15000 $Y=16500 $D=1
M3 10 4 12 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=15000 $Y=32700 $D=1
M4 39 en 10 10 n L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=21600 $Y=16500 $D=1
M5 19 12 10 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=21600 $Y=29700 $D=1
M6 14 clk 39 10 n L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=23100 $Y=16500 $D=1
M7 10 fa_in 19 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=24000 $Y=29700 $D=1
M8 40 14 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=28800 $Y=19500 $D=1
M9 16 13 19 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=4.5e-12 PD=9e-06 PS=9e-06 $X=28800 $Y=29700 $D=1
M10 15 14 40 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=30300 $Y=19500 $D=1
M11 41 fa_in 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=33600 $Y=29700 $D=1
M12 42 11 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=35100 $Y=19500 $D=1
M13 16 12 41 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=35100 $Y=29700 $D=1
M14 21 14 42 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=2.7e-12 PD=9.6e-06 PS=7.8e-06 $X=36600 $Y=19500 $D=1
M15 43 15 21 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=5.4e-12 PD=7.8e-06 PS=9.6e-06 $X=39000 $Y=19500 $D=1
M16 23 13 10 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=39900 $Y=29700 $D=1
M17 10 22 43 10 n L=6e-07 W=3e-06 AD=6.3e-12 AS=2.7e-12 PD=1.02e-05 PS=7.8e-06 $X=40500 $Y=19500 $D=1
M18 10 fa_in 23 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=5.4e-12 PD=9.6e-06 PS=9.6e-06 $X=42300 $Y=29700 $D=1
M19 22 21 10 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=6.3e-12 PD=9e-06 PS=1.02e-05 $X=43200 $Y=19500 $D=1
M20 23 12 10 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=44700 $Y=29700 $D=1
M21 44 22 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=48000 $Y=19500 $D=1
M22 25 15 44 10 n L=6e-07 W=3e-06 AD=5.4e-12 AS=2.7e-12 PD=9.6e-06 PS=7.8e-06 $X=49500 $Y=19500 $D=1
M23 27 16 23 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=4.5e-12 PD=9e-06 PS=9e-06 $X=49500 $Y=29700 $D=1
M24 45 14 25 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=5.4e-12 PD=7.8e-06 PS=9.6e-06 $X=51900 $Y=19500 $D=1
M25 10 Out 45 10 n L=6e-07 W=3e-06 AD=6.3e-12 AS=2.7e-12 PD=1.02e-05 PS=7.8e-06 $X=53400 $Y=19500 $D=1
M26 46 13 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=4.5e-12 PD=7.8e-06 PS=9e-06 $X=54300 $Y=29700 $D=1
M27 47 fa_in 46 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=2.7e-12 PD=7.8e-06 PS=7.8e-06 $X=55800 $Y=29700 $D=1
M28 48 25 10 10 n L=6e-07 W=3e-06 AD=2.7e-12 AS=6.3e-12 PD=7.8e-06 PS=1.02e-05 $X=56100 $Y=19500 $D=1
M29 27 12 47 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=57300 $Y=29700 $D=1
M30 Out 25 48 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=2.7e-12 PD=9e-06 PS=7.8e-06 $X=57600 $Y=19500 $D=1
M31 17 27 10 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=4.5e-12 PD=9e-06 PS=9e-06 $X=62100 $Y=29700 $D=1
M32 Cout 16 10 10 n L=6e-07 W=3e-06 AD=4.5e-12 AS=4.5e-12 PD=9e-06 PS=9e-06 $X=66900 $Y=29700 $D=1
M33 11 4 5 26 p L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=12600 $Y=3900 $D=0
M34 12 4 6 Cin p L=6e-07 W=3e-06 AD=5.4e-12 AS=4.5e-12 PD=9.6e-06 PS=9e-06 $X=12600 $Y=45300 $D=0
M35 3 8 11 26 p L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=15000 $Y=3900 $D=0
M36 10 9 12 Cin p L=6e-07 W=3e-06 AD=4.5e-12 AS=5.4e-12 PD=9e-06 PS=9.6e-06 $X=15000 $Y=45300 $D=0
M37 14 en 26 26 p L=6e-07 W=6e-06 AD=1.08e-11 AS=9e-12 PD=1.56e-05 PS=1.5e-05 $X=21600 $Y=2700 $D=0
M38 20 12 Cin Cin p L=6e-07 W=6e-06 AD=1.08e-11 AS=9e-12 PD=1.56e-05 PS=1.5e-05 $X=21600 $Y=43500 $D=0
M39 26 clk 14 26 p L=6e-07 W=6e-06 AD=9e-12 AS=1.08e-11 PD=1.5e-05 PS=1.56e-05 $X=24000 $Y=2700 $D=0
M40 Cin fa_in 20 Cin p L=6e-07 W=6e-06 AD=9e-12 AS=1.08e-11 PD=1.5e-05 PS=1.56e-05 $X=24000 $Y=43500 $D=0
M41 30 14 26 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=28800 $Y=2700 $D=0
M42 16 13 20 Cin p L=6e-07 W=6e-06 AD=9e-12 AS=9e-12 PD=1.5e-05 PS=1.5e-05 $X=28800 $Y=43500 $D=0
M43 15 14 30 26 p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=30300 $Y=2700 $D=0
M44 31 fa_in Cin Cin p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=33600 $Y=43500 $D=0
M45 32 11 26 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=35100 $Y=2700 $D=0
M46 16 12 31 Cin p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=35100 $Y=43500 $D=0
M47 21 15 32 26 p L=6e-07 W=6e-06 AD=1.08e-11 AS=5.4e-12 PD=1.56e-05 PS=1.38e-05 $X=36600 $Y=2700 $D=0
M48 33 14 21 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.08e-11 PD=1.38e-05 PS=1.56e-05 $X=39000 $Y=2700 $D=0
M49 24 13 Cin Cin p L=6e-07 W=6e-06 AD=1.08e-11 AS=9e-12 PD=1.56e-05 PS=1.5e-05 $X=39900 $Y=43500 $D=0
M50 26 22 33 26 p L=6e-07 W=6e-06 AD=1.26e-11 AS=5.4e-12 PD=1.62e-05 PS=1.38e-05 $X=40500 $Y=2700 $D=0
M51 Cin fa_in 24 Cin p L=6e-07 W=6e-06 AD=1.08e-11 AS=1.08e-11 PD=1.56e-05 PS=1.56e-05 $X=42300 $Y=43500 $D=0
M52 22 21 26 26 p L=6e-07 W=6e-06 AD=9e-12 AS=1.26e-11 PD=1.5e-05 PS=1.62e-05 $X=43200 $Y=2700 $D=0
M53 24 12 Cin Cin p L=6e-07 W=6e-06 AD=9e-12 AS=1.08e-11 PD=1.5e-05 PS=1.56e-05 $X=44700 $Y=43500 $D=0
M54 34 22 26 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=48000 $Y=2700 $D=0
M55 25 14 34 26 p L=6e-07 W=6e-06 AD=1.08e-11 AS=5.4e-12 PD=1.56e-05 PS=1.38e-05 $X=49500 $Y=2700 $D=0
M56 27 16 24 Cin p L=6e-07 W=6e-06 AD=9e-12 AS=9e-12 PD=1.5e-05 PS=1.5e-05 $X=49500 $Y=43500 $D=0
M57 35 15 25 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.08e-11 PD=1.38e-05 PS=1.56e-05 $X=51900 $Y=2700 $D=0
M58 26 Out 35 26 p L=6e-07 W=6e-06 AD=1.26e-11 AS=5.4e-12 PD=1.62e-05 PS=1.38e-05 $X=53400 $Y=2700 $D=0
M59 36 13 Cin Cin p L=6e-07 W=6e-06 AD=5.4e-12 AS=9e-12 PD=1.38e-05 PS=1.5e-05 $X=54300 $Y=43500 $D=0
M60 37 fa_in 36 Cin p L=6e-07 W=6e-06 AD=5.4e-12 AS=5.4e-12 PD=1.38e-05 PS=1.38e-05 $X=55800 $Y=43500 $D=0
M61 38 25 26 26 p L=6e-07 W=6e-06 AD=5.4e-12 AS=1.26e-11 PD=1.38e-05 PS=1.62e-05 $X=56100 $Y=2700 $D=0
M62 27 12 37 Cin p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=57300 $Y=43500 $D=0
M63 Out 25 38 26 p L=6e-07 W=6e-06 AD=9e-12 AS=5.4e-12 PD=1.5e-05 PS=1.38e-05 $X=57600 $Y=2700 $D=0
M64 17 27 Cin Cin p L=6e-07 W=6e-06 AD=9e-12 AS=9e-12 PD=1.5e-05 PS=1.5e-05 $X=62100 $Y=43500 $D=0
M65 Cout 16 Cin Cin p L=6e-07 W=6e-06 AD=9e-12 AS=9e-12 PD=1.5e-05 PS=1.5e-05 $X=66900 $Y=43500 $D=0
X66 4 10 26 8 ______inv_magic_inverter $T=3900 24900 1 0 $X=2400 $Y=-600
X67 4 10 Cin 9 ______inv_magic_inverter $T=3900 27300 0 0 $X=2400 $Y=26400
.ENDS
***************************************
