magic
tech scmos
timestamp 1543271335
<< metal1 >>
rect -1 174 244 177
rect 64 168 69 174
rect 236 168 244 174
rect -1 145 8 149
rect 64 83 244 96
rect 64 78 87 83
rect 93 78 244 83
rect 86 54 87 58
rect 73 48 74 52
rect 199 42 244 47
rect -1 24 8 28
rect -1 17 8 21
rect -1 1 87 6
rect 93 1 244 6
rect -1 -3 244 1
<< m2contact >>
rect 8 145 12 149
rect 74 48 78 52
rect 67 38 71 42
rect 8 24 12 28
rect 8 17 12 21
<< metal2 >>
rect 12 145 79 149
rect 75 123 79 145
rect 75 119 88 123
rect 60 112 67 116
rect 60 102 64 112
rect 64 71 87 75
rect 67 28 71 38
rect 12 24 71 28
rect 74 21 78 48
rect 12 17 78 21
use ../../fa/magic/fa  fa_0 ../../fa/magic
timestamp 1542251572
transform 1 0 61 0 1 90
box 0 -4 175 89
use ../../bc1a/magic/bc1a  bc1a_0 ../../bc1a/magic
timestamp 1542169151
transform 1 0 0 0 1 12
box -1 -12 64 162
use ../../nand/magic/nand  nand_0 ../../nand/magic
timestamp 1543271335
transform 1 0 65 0 -1 81
box -4 -3 28 81
use ../../dffpos/magic/dffpos  dffpos_0 ../../dffpos/magic
timestamp 1543271063
transform 1 0 63 0 1 0
box 18 0 139 84
<< labels >>
rlabel metal1 176 176 176 176 5 c_in
rlabel metal1 1 147 1 147 3 fa_in
rlabel metal1 1 26 1 26 3 clk
rlabel metal1 1 19 1 19 3 en
<< end >>
