magic
tech scmos
timestamp 1542725905
<< metal1 >>
rect -24 22 24 24
rect -24 -22 -22 22
rect 22 -22 24 22
rect -24 -24 24 -22
<< m2contact >>
rect -22 -22 22 22
<< metal2 >>
rect -24 22 24 24
rect -24 -22 -22 22
rect 22 -22 24 22
rect -24 -24 24 -22
<< end >>
